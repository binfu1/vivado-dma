`timescale 1ns / 1ns
`define SYNTH
//////////////////////////////////////////////////////////////////////////////////
// Company: 浪潮信息
// Engineer: 邓子为
//////////////////////////////////////////////////////////////////////////////////

module top #(
  parameter SIZE_LOOP = 128  //计算的平面数量
  ) (
`ifdef SYNTH
  input         init_clk,      //初始化时钟
  input         sys_clk_clk_p, //PCIe时钟
  input         sys_clk_clk_n,
  input         sys_rstn,      //PCIe复位
  input  [15:0] pcie_mgt_rxn,  //PCIe引脚
  input  [15:0] pcie_mgt_rxp,
  output [15:0] pcie_mgt_txn,
  output [15:0] pcie_mgt_txp
`else
  input         sclk,  
  input         xdma_rstn, 
  input  [31:0] gpio
`endif
);

localparam LENGTH      = 128; //FFT的点数
localparam FFT_NUM     = 8;  //FFT核数量
localparam DWIDTH_FFT  = 32; //FFT数据实部和虚部位宽，BIT
localparam DWIDTH_BRAM = 64; //本地内存的数据位宽，BIT
localparam AWIDTH_BRAM = 14; //本地内存的地址位宽
localparam AWIDTH_HBM  = 32; //全局内存的地址位宽
localparam DWIDTH_HBM  = 32; //全局内存的数据位宽，BYTE
localparam NUM_GROUP   = 16;  //分组数量
localparam SIZE_GROUP  = LENGTH/NUM_GROUP;

/**************************** XDMA系统 ****************************/
wire    [NUM_GROUP-1:0] m_axi_awready;
wire    [NUM_GROUP-1:0] m_axi_awvalid;
wire   [AWIDTH_HBM-1:0] m_axi_awaddr  [NUM_GROUP-1:0];
wire              [1:0] m_axi_awburst [NUM_GROUP-1:0];
wire              [3:0] m_axi_awcache [NUM_GROUP-1:0];
wire              [7:0] m_axi_awlen   [NUM_GROUP-1:0];
wire              [2:0] m_axi_awsize  [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] m_axi_wready;
wire    [NUM_GROUP-1:0] m_axi_wvalid;
wire [DWIDTH_HBM*8-1:0] m_axi_wdata   [NUM_GROUP-1:0];
wire   [DWIDTH_HBM-1:0] m_axi_wstrb   [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] m_axi_wlast;
wire    [NUM_GROUP-1:0] m_axi_bready;
wire    [NUM_GROUP-1:0] m_axi_bvalid;
wire              [1:0] m_axi_bresp   [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] m_axi_arready;
wire    [NUM_GROUP-1:0] m_axi_arvalid;
wire   [AWIDTH_HBM-1:0] m_axi_araddr  [NUM_GROUP-1:0];
wire              [1:0] m_axi_arburst [NUM_GROUP-1:0];
wire              [3:0] m_axi_arcache [NUM_GROUP-1:0];
wire              [7:0] m_axi_arlen   [NUM_GROUP-1:0];
wire              [2:0] m_axi_arsize  [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] m_axi_rready;
wire    [NUM_GROUP-1:0] m_axi_rvalid;
wire [DWIDTH_HBM*8-1:0] m_axi_rdata   [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] m_axi_rlast;
wire              [1:0] m_axi_rresp   [NUM_GROUP-1:0];

`ifdef SYNTH
wire [31:0] gpio;
xdma_wrapper xdma_wrapper_i(
  .hbm_refclk     (init_clk),
  .pcie_mgt_rxn   (pcie_mgt_rxn),
  .pcie_mgt_rxp   (pcie_mgt_rxp),
  .pcie_mgt_txn   (pcie_mgt_txn),
  .pcie_mgt_txp   (pcie_mgt_txp),
  .sys_clk_clk_n  (sys_clk_clk_n),
  .sys_clk_clk_p  (sys_clk_clk_p),
  .sys_rstn       (sys_rstn),
  .xdma_aclk      (sclk),
  .xdma_rstn      (xdma_rstn),
  .gpio           (gpio), 
  .msi_enable     (msi_enable),
  .irq_req        (irq_req),

  .cu_axi0_awready (m_axi_awready[0]),
  .cu_axi0_awvalid (m_axi_awvalid[0]),
  .cu_axi0_awaddr  (m_axi_awaddr [0]),
  .cu_axi0_wready  (m_axi_wready [0]),
  .cu_axi0_wvalid  (m_axi_wvalid [0]),
  .cu_axi0_wdata   (m_axi_wdata  [0]),
  .cu_axi0_wstrb   (m_axi_wstrb  [0]),
  .cu_axi0_wlast   (m_axi_wlast  [0]),
  .cu_axi0_bready  (m_axi_bready [0]),
  .cu_axi0_bvalid  (m_axi_bvalid [0]),
  .cu_axi0_bresp   (m_axi_bresp  [0]),
  .cu_axi0_awburst (m_axi_awburst[0]),
  .cu_axi0_awcache (m_axi_awcache[0]),
  .cu_axi0_awlen   (m_axi_awlen  [0]),
  .cu_axi0_awsize  (m_axi_awsize [0]),
  .cu_axi0_arready (m_axi_arready[0]),
  .cu_axi0_arvalid (m_axi_arvalid[0]),
  .cu_axi0_araddr  (m_axi_araddr [0]),
  .cu_axi0_rready  (m_axi_rready [0]),
  .cu_axi0_rvalid  (m_axi_rvalid [0]),
  .cu_axi0_rdata   (m_axi_rdata  [0]),
  .cu_axi0_rlast   (m_axi_rlast  [0]),
  .cu_axi0_rresp   (m_axi_rresp  [0]),
  .cu_axi0_arburst (m_axi_arburst[0]),
  .cu_axi0_arcache (m_axi_arcache[0]),
  .cu_axi0_arlen   (m_axi_arlen  [0]),
  .cu_axi0_arsize  (m_axi_arsize [0]),
  //.cu_axi0_awid    (),
  .cu_axi0_awprot  (),
  .cu_axi0_awlock  (),
  .cu_axi0_awqos   (),
  .cu_axi0_awregion(),
  //.cu_axi0_arid    (),
  .cu_axi0_arprot  (),
  .cu_axi0_arlock  (),
  .cu_axi0_arqos   (),
  .cu_axi0_arregion(),
  //.cu_axi0_bid     (),
  //.cu_axi0_rid     (),

  .cu_axi1_awready (m_axi_awready[1]),
  .cu_axi1_awvalid (m_axi_awvalid[1]),
  .cu_axi1_awaddr  (m_axi_awaddr [1]),
  .cu_axi1_wready  (m_axi_wready [1]),
  .cu_axi1_wvalid  (m_axi_wvalid [1]),
  .cu_axi1_wdata   (m_axi_wdata  [1]),
  .cu_axi1_wstrb   (m_axi_wstrb  [1]),
  .cu_axi1_wlast   (m_axi_wlast  [1]),
  .cu_axi1_bready  (m_axi_bready [1]),
  .cu_axi1_bvalid  (m_axi_bvalid [1]),
  .cu_axi1_bresp   (m_axi_bresp  [1]),
  .cu_axi1_awburst (m_axi_awburst[1]),
  .cu_axi1_awcache (m_axi_awcache[1]),
  .cu_axi1_awlen   (m_axi_awlen  [1]),
  .cu_axi1_awsize  (m_axi_awsize [1]),
  .cu_axi1_arready (m_axi_arready[1]),
  .cu_axi1_arvalid (m_axi_arvalid[1]),
  .cu_axi1_araddr  (m_axi_araddr [1]),
  .cu_axi1_rready  (m_axi_rready [1]),
  .cu_axi1_rvalid  (m_axi_rvalid [1]),
  .cu_axi1_rdata   (m_axi_rdata  [1]),
  .cu_axi1_rlast   (m_axi_rlast  [1]),
  .cu_axi1_rresp   (m_axi_rresp  [1]),
  .cu_axi1_arburst (m_axi_arburst[1]),
  .cu_axi1_arcache (m_axi_arcache[1]),
  .cu_axi1_arlen   (m_axi_arlen  [1]),
  .cu_axi1_arsize  (m_axi_arsize [1]),
  //.cu_axi1_awid    (),
  .cu_axi1_awprot  (),
  .cu_axi1_awlock  (),
  .cu_axi1_awqos   (),
  .cu_axi1_awregion(),
  //.cu_axi1_arid    (),
  .cu_axi1_arprot  (),
  .cu_axi1_arlock  (),
  .cu_axi1_arqos   (),
  .cu_axi1_arregion(),
  //.cu_axi1_bid     (),
  //.cu_axi1_rid     (),

  .cu_axi2_awready (m_axi_awready[2]),
  .cu_axi2_awvalid (m_axi_awvalid[2]),
  .cu_axi2_awaddr  (m_axi_awaddr [2]),
  .cu_axi2_wready  (m_axi_wready [2]),
  .cu_axi2_wvalid  (m_axi_wvalid [2]),
  .cu_axi2_wdata   (m_axi_wdata  [2]),
  .cu_axi2_wstrb   (m_axi_wstrb  [2]),
  .cu_axi2_wlast   (m_axi_wlast  [2]),
  .cu_axi2_bready  (m_axi_bready [2]),
  .cu_axi2_bvalid  (m_axi_bvalid [2]),
  .cu_axi2_bresp   (m_axi_bresp  [2]),
  .cu_axi2_awburst (m_axi_awburst[2]),
  .cu_axi2_awcache (m_axi_awcache[2]),
  .cu_axi2_awlen   (m_axi_awlen  [2]),
  .cu_axi2_awsize  (m_axi_awsize [2]),
  .cu_axi2_arready (m_axi_arready[2]),
  .cu_axi2_arvalid (m_axi_arvalid[2]),
  .cu_axi2_araddr  (m_axi_araddr [2]),
  .cu_axi2_rready  (m_axi_rready [2]),
  .cu_axi2_rvalid  (m_axi_rvalid [2]),
  .cu_axi2_rdata   (m_axi_rdata  [2]),
  .cu_axi2_rlast   (m_axi_rlast  [2]),
  .cu_axi2_rresp   (m_axi_rresp  [2]),
  .cu_axi2_arburst (m_axi_arburst[2]),
  .cu_axi2_arcache (m_axi_arcache[2]),
  .cu_axi2_arlen   (m_axi_arlen  [2]),
  .cu_axi2_arsize  (m_axi_arsize [2]),
  //.cu_axi2_awid    (),
  .cu_axi2_awprot  (),
  .cu_axi2_awlock  (),
  .cu_axi2_awqos   (),
  .cu_axi2_awregion(),
  //.cu_axi2_arid    (),
  .cu_axi2_arprot  (),
  .cu_axi2_arlock  (),
  .cu_axi2_arqos   (),
  .cu_axi2_arregion(),
  //.cu_axi2_bid     (),
  //.cu_axi2_rid     (),

  .cu_axi3_awready (m_axi_awready[3]),
  .cu_axi3_awvalid (m_axi_awvalid[3]),
  .cu_axi3_awaddr  (m_axi_awaddr [3]),
  .cu_axi3_wready  (m_axi_wready [3]),
  .cu_axi3_wvalid  (m_axi_wvalid [3]),
  .cu_axi3_wdata   (m_axi_wdata  [3]),
  .cu_axi3_wstrb   (m_axi_wstrb  [3]),
  .cu_axi3_wlast   (m_axi_wlast  [3]),
  .cu_axi3_bready  (m_axi_bready [3]),
  .cu_axi3_bvalid  (m_axi_bvalid [3]),
  .cu_axi3_bresp   (m_axi_bresp  [3]),
  .cu_axi3_awburst (m_axi_awburst[3]),
  .cu_axi3_awcache (m_axi_awcache[3]),
  .cu_axi3_awlen   (m_axi_awlen  [3]),
  .cu_axi3_awsize  (m_axi_awsize [3]),
  .cu_axi3_arready (m_axi_arready[3]),
  .cu_axi3_arvalid (m_axi_arvalid[3]),
  .cu_axi3_araddr  (m_axi_araddr [3]),
  .cu_axi3_rready  (m_axi_rready [3]),
  .cu_axi3_rvalid  (m_axi_rvalid [3]),
  .cu_axi3_rdata   (m_axi_rdata  [3]),
  .cu_axi3_rlast   (m_axi_rlast  [3]),
  .cu_axi3_rresp   (m_axi_rresp  [3]),
  .cu_axi3_arburst (m_axi_arburst[3]),
  .cu_axi3_arcache (m_axi_arcache[3]),
  .cu_axi3_arlen   (m_axi_arlen  [3]),
  .cu_axi3_arsize  (m_axi_arsize [3]),
  //.cu_axi3_awid    (),
  .cu_axi3_awprot  (),
  .cu_axi3_awlock  (),
  .cu_axi3_awqos   (),
  .cu_axi3_awregion(),
  //.cu_axi3_arid    (),
  .cu_axi3_arprot  (),
  .cu_axi3_arlock  (),
  .cu_axi3_arqos   (),
  .cu_axi3_arregion(),
  //.cu_axi3_bid     (),
  //.cu_axi3_rid     (),

  .cu_axi4_awready (m_axi_awready[4]),
  .cu_axi4_awvalid (m_axi_awvalid[4]),
  .cu_axi4_awaddr  (m_axi_awaddr [4]),
  .cu_axi4_wready  (m_axi_wready [4]),
  .cu_axi4_wvalid  (m_axi_wvalid [4]),
  .cu_axi4_wdata   (m_axi_wdata  [4]),
  .cu_axi4_wstrb   (m_axi_wstrb  [4]),
  .cu_axi4_wlast   (m_axi_wlast  [4]),
  .cu_axi4_bready  (m_axi_bready [4]),
  .cu_axi4_bvalid  (m_axi_bvalid [4]),
  .cu_axi4_bresp   (m_axi_bresp  [4]),
  .cu_axi4_awburst (m_axi_awburst[4]),
  .cu_axi4_awcache (m_axi_awcache[4]),
  .cu_axi4_awlen   (m_axi_awlen  [4]),
  .cu_axi4_awsize  (m_axi_awsize [4]),
  .cu_axi4_arready (m_axi_arready[4]),
  .cu_axi4_arvalid (m_axi_arvalid[4]),
  .cu_axi4_araddr  (m_axi_araddr [4]),
  .cu_axi4_rready  (m_axi_rready [4]),
  .cu_axi4_rvalid  (m_axi_rvalid [4]),
  .cu_axi4_rdata   (m_axi_rdata  [4]),
  .cu_axi4_rlast   (m_axi_rlast  [4]),
  .cu_axi4_rresp   (m_axi_rresp  [4]),
  .cu_axi4_arburst (m_axi_arburst[4]),
  .cu_axi4_arcache (m_axi_arcache[4]),
  .cu_axi4_arlen   (m_axi_arlen  [4]),
  .cu_axi4_arsize  (m_axi_arsize [4]),
  //.cu_axi4_awid    (),
  .cu_axi4_awprot  (),
  .cu_axi4_awlock  (),
  .cu_axi4_awqos   (),
  .cu_axi4_awregion(),
  //.cu_axi4_arid    (),
  .cu_axi4_arprot  (),
  .cu_axi4_arlock  (),
  .cu_axi4_arqos   (),
  .cu_axi4_arregion(),
  //.cu_axi4_bid     (),
  //.cu_axi4_rid     (),

  .cu_axi5_awready (m_axi_awready[5]),
  .cu_axi5_awvalid (m_axi_awvalid[5]),
  .cu_axi5_awaddr  (m_axi_awaddr [5]),
  .cu_axi5_wready  (m_axi_wready [5]),
  .cu_axi5_wvalid  (m_axi_wvalid [5]),
  .cu_axi5_wdata   (m_axi_wdata  [5]),
  .cu_axi5_wstrb   (m_axi_wstrb  [5]),
  .cu_axi5_wlast   (m_axi_wlast  [5]),
  .cu_axi5_bready  (m_axi_bready [5]),
  .cu_axi5_bvalid  (m_axi_bvalid [5]),
  .cu_axi5_bresp   (m_axi_bresp  [5]),
  .cu_axi5_awburst (m_axi_awburst[5]),
  .cu_axi5_awcache (m_axi_awcache[5]),
  .cu_axi5_awlen   (m_axi_awlen  [5]),
  .cu_axi5_awsize  (m_axi_awsize [5]),
  .cu_axi5_arready (m_axi_arready[5]),
  .cu_axi5_arvalid (m_axi_arvalid[5]),
  .cu_axi5_araddr  (m_axi_araddr [5]),
  .cu_axi5_rready  (m_axi_rready [5]),
  .cu_axi5_rvalid  (m_axi_rvalid [5]),
  .cu_axi5_rdata   (m_axi_rdata  [5]),
  .cu_axi5_rlast   (m_axi_rlast  [5]),
  .cu_axi5_rresp   (m_axi_rresp  [5]),
  .cu_axi5_arburst (m_axi_arburst[5]),
  .cu_axi5_arcache (m_axi_arcache[5]),
  .cu_axi5_arlen   (m_axi_arlen  [5]),
  .cu_axi5_arsize  (m_axi_arsize [5]),
  //.cu_axi5_awid    (),
  .cu_axi5_awprot  (),
  .cu_axi5_awlock  (),
  .cu_axi5_awqos   (),
  .cu_axi5_awregion(),
  //.cu_axi5_arid    (),
  .cu_axi5_arprot  (),
  .cu_axi5_arlock  (),
  .cu_axi5_arqos   (),
  .cu_axi5_arregion(),
  //.cu_axi5_bid     (),
  //.cu_axi5_rid     (),

  .cu_axi6_awready (m_axi_awready[6]),
  .cu_axi6_awvalid (m_axi_awvalid[6]),
  .cu_axi6_awaddr  (m_axi_awaddr [6]),
  .cu_axi6_wready  (m_axi_wready [6]),
  .cu_axi6_wvalid  (m_axi_wvalid [6]),
  .cu_axi6_wdata   (m_axi_wdata  [6]),
  .cu_axi6_wstrb   (m_axi_wstrb  [6]),
  .cu_axi6_wlast   (m_axi_wlast  [6]),
  .cu_axi6_bready  (m_axi_bready [6]),
  .cu_axi6_bvalid  (m_axi_bvalid [6]),
  .cu_axi6_bresp   (m_axi_bresp  [6]),
  .cu_axi6_awburst (m_axi_awburst[6]),
  .cu_axi6_awcache (m_axi_awcache[6]),
  .cu_axi6_awlen   (m_axi_awlen  [6]),
  .cu_axi6_awsize  (m_axi_awsize [6]),
  .cu_axi6_arready (m_axi_arready[6]),
  .cu_axi6_arvalid (m_axi_arvalid[6]),
  .cu_axi6_araddr  (m_axi_araddr [6]),
  .cu_axi6_rready  (m_axi_rready [6]),
  .cu_axi6_rvalid  (m_axi_rvalid [6]),
  .cu_axi6_rdata   (m_axi_rdata  [6]),
  .cu_axi6_rlast   (m_axi_rlast  [6]),
  .cu_axi6_rresp   (m_axi_rresp  [6]),
  .cu_axi6_arburst (m_axi_arburst[6]),
  .cu_axi6_arcache (m_axi_arcache[6]),
  .cu_axi6_arlen   (m_axi_arlen  [6]),
  .cu_axi6_arsize  (m_axi_arsize [6]),
  //.cu_axi6_awid    (),
  .cu_axi6_awprot  (),
  .cu_axi6_awlock  (),
  .cu_axi6_awqos   (),
  .cu_axi6_awregion(),
  //.cu_axi6_arid    (),
  .cu_axi6_arprot  (),
  .cu_axi6_arlock  (),
  .cu_axi6_arqos   (),
  .cu_axi6_arregion(),
  //.cu_axi6_bid     (),
  //.cu_axi6_rid     (),

  .cu_axi7_awready (m_axi_awready[7]),
  .cu_axi7_awvalid (m_axi_awvalid[7]),
  .cu_axi7_awaddr  (m_axi_awaddr [7]),
  .cu_axi7_wready  (m_axi_wready [7]),
  .cu_axi7_wvalid  (m_axi_wvalid [7]),
  .cu_axi7_wdata   (m_axi_wdata  [7]),
  .cu_axi7_wstrb   (m_axi_wstrb  [7]),
  .cu_axi7_wlast   (m_axi_wlast  [7]),
  .cu_axi7_bready  (m_axi_bready [7]),
  .cu_axi7_bvalid  (m_axi_bvalid [7]),
  .cu_axi7_bresp   (m_axi_bresp  [7]),
  .cu_axi7_awburst (m_axi_awburst[7]),
  .cu_axi7_awcache (m_axi_awcache[7]),
  .cu_axi7_awlen   (m_axi_awlen  [7]),
  .cu_axi7_awsize  (m_axi_awsize [7]),
  .cu_axi7_arready (m_axi_arready[7]),
  .cu_axi7_arvalid (m_axi_arvalid[7]),
  .cu_axi7_araddr  (m_axi_araddr [7]),
  .cu_axi7_rready  (m_axi_rready [7]),
  .cu_axi7_rvalid  (m_axi_rvalid [7]),
  .cu_axi7_rdata   (m_axi_rdata  [7]),
  .cu_axi7_rlast   (m_axi_rlast  [7]),
  .cu_axi7_rresp   (m_axi_rresp  [7]),
  .cu_axi7_arburst (m_axi_arburst[7]),
  .cu_axi7_arcache (m_axi_arcache[7]),
  .cu_axi7_arlen   (m_axi_arlen  [7]),
  .cu_axi7_arsize  (m_axi_arsize [7]),
  //.cu_axi7_awid    (),
  .cu_axi7_awprot  (),
  .cu_axi7_awlock  (),
  .cu_axi7_awqos   (),
  .cu_axi7_awregion(),
  //.cu_axi7_arid    (),
  .cu_axi7_arprot  (),
  .cu_axi7_arlock  (),
  .cu_axi7_arqos   (),
  .cu_axi7_arregion(),
  //.cu_axi7_bid     (),
  //.cu_axi7_rid     (),

  .cu_axi8_awready (m_axi_awready[8]),
  .cu_axi8_awvalid (m_axi_awvalid[8]),
  .cu_axi8_awaddr  (m_axi_awaddr [8]),
  .cu_axi8_wready  (m_axi_wready [8]),
  .cu_axi8_wvalid  (m_axi_wvalid [8]),
  .cu_axi8_wdata   (m_axi_wdata  [8]),
  .cu_axi8_wstrb   (m_axi_wstrb  [8]),
  .cu_axi8_wlast   (m_axi_wlast  [8]),
  .cu_axi8_bready  (m_axi_bready [8]),
  .cu_axi8_bvalid  (m_axi_bvalid [8]),
  .cu_axi8_bresp   (m_axi_bresp  [8]),
  .cu_axi8_awburst (m_axi_awburst[8]),
  .cu_axi8_awcache (m_axi_awcache[8]),
  .cu_axi8_awlen   (m_axi_awlen  [8]),
  .cu_axi8_awsize  (m_axi_awsize [8]),
  .cu_axi8_arready (m_axi_arready[8]),
  .cu_axi8_arvalid (m_axi_arvalid[8]),
  .cu_axi8_araddr  (m_axi_araddr [8]),
  .cu_axi8_rready  (m_axi_rready [8]),
  .cu_axi8_rvalid  (m_axi_rvalid [8]),
  .cu_axi8_rdata   (m_axi_rdata  [8]),
  .cu_axi8_rlast   (m_axi_rlast  [8]),
  .cu_axi8_rresp   (m_axi_rresp  [8]),
  .cu_axi8_arburst (m_axi_arburst[8]),
  .cu_axi8_arcache (m_axi_arcache[8]),
  .cu_axi8_arlen   (m_axi_arlen  [8]),
  .cu_axi8_arsize  (m_axi_arsize [8]),
  //.cu_axi8_awid    (),
  .cu_axi8_awprot  (),
  .cu_axi8_awlock  (),
  .cu_axi8_awqos   (),
  .cu_axi8_awregion(),
  //.cu_axi8_arid    (),
  .cu_axi8_arprot  (),
  .cu_axi8_arlock  (),
  .cu_axi8_arqos   (),
  .cu_axi8_arregion(),
  //.cu_axi8_bid     (),
  //.cu_axi8_rid     (),

  .cu_axi9_awready (m_axi_awready[9]),
  .cu_axi9_awvalid (m_axi_awvalid[9]),
  .cu_axi9_awaddr  (m_axi_awaddr [9]),
  .cu_axi9_wready  (m_axi_wready [9]),
  .cu_axi9_wvalid  (m_axi_wvalid [9]),
  .cu_axi9_wdata   (m_axi_wdata  [9]),
  .cu_axi9_wstrb   (m_axi_wstrb  [9]),
  .cu_axi9_wlast   (m_axi_wlast  [9]),
  .cu_axi9_bready  (m_axi_bready [9]),
  .cu_axi9_bvalid  (m_axi_bvalid [9]),
  .cu_axi9_bresp   (m_axi_bresp  [9]),
  .cu_axi9_awburst (m_axi_awburst[9]),
  .cu_axi9_awcache (m_axi_awcache[9]),
  .cu_axi9_awlen   (m_axi_awlen  [9]),
  .cu_axi9_awsize  (m_axi_awsize [9]),
  .cu_axi9_arready (m_axi_arready[9]),
  .cu_axi9_arvalid (m_axi_arvalid[9]),
  .cu_axi9_araddr  (m_axi_araddr [9]),
  .cu_axi9_rready  (m_axi_rready [9]),
  .cu_axi9_rvalid  (m_axi_rvalid [9]),
  .cu_axi9_rdata   (m_axi_rdata  [9]),
  .cu_axi9_rlast   (m_axi_rlast  [9]),
  .cu_axi9_rresp   (m_axi_rresp  [9]),
  .cu_axi9_arburst (m_axi_arburst[9]),
  .cu_axi9_arcache (m_axi_arcache[9]),
  .cu_axi9_arlen   (m_axi_arlen  [9]),
  .cu_axi9_arsize  (m_axi_arsize [9]),
  //.cu_axi9_awid    (),
  .cu_axi9_awprot  (),
  .cu_axi9_awlock  (),
  .cu_axi9_awqos   (),
  .cu_axi9_awregion(),
  //.cu_axi9_arid    (),
  .cu_axi9_arprot  (),
  .cu_axi9_arlock  (),
  .cu_axi9_arqos   (),
  .cu_axi9_arregion(),
  //.cu_axi9_bid     (),
  //.cu_axi9_rid     (),

  .cu_axi10_awready (m_axi_awready[10]),
  .cu_axi10_awvalid (m_axi_awvalid[10]),
  .cu_axi10_awaddr  (m_axi_awaddr [10]),
  .cu_axi10_wready  (m_axi_wready [10]),
  .cu_axi10_wvalid  (m_axi_wvalid [10]),
  .cu_axi10_wdata   (m_axi_wdata  [10]),
  .cu_axi10_wstrb   (m_axi_wstrb  [10]),
  .cu_axi10_wlast   (m_axi_wlast  [10]),
  .cu_axi10_bready  (m_axi_bready [10]),
  .cu_axi10_bvalid  (m_axi_bvalid [10]),
  .cu_axi10_bresp   (m_axi_bresp  [10]),
  .cu_axi10_awburst (m_axi_awburst[10]),
  .cu_axi10_awcache (m_axi_awcache[10]),
  .cu_axi10_awlen   (m_axi_awlen  [10]),
  .cu_axi10_awsize  (m_axi_awsize [10]),
  .cu_axi10_arready (m_axi_arready[10]),
  .cu_axi10_arvalid (m_axi_arvalid[10]),
  .cu_axi10_araddr  (m_axi_araddr [10]),
  .cu_axi10_rready  (m_axi_rready [10]),
  .cu_axi10_rvalid  (m_axi_rvalid [10]),
  .cu_axi10_rdata   (m_axi_rdata  [10]),
  .cu_axi10_rlast   (m_axi_rlast  [10]),
  .cu_axi10_rresp   (m_axi_rresp  [10]),
  .cu_axi10_arburst (m_axi_arburst[10]),
  .cu_axi10_arcache (m_axi_arcache[10]),
  .cu_axi10_arlen   (m_axi_arlen  [10]),
  .cu_axi10_arsize  (m_axi_arsize [10]),
  //.cu_axi10_awid    (),
  .cu_axi10_awprot  (),
  .cu_axi10_awlock  (),
  .cu_axi10_awqos   (),
  .cu_axi10_awregion(),
  //.cu_axi10_arid    (),
  .cu_axi10_arprot  (),
  .cu_axi10_arlock  (),
  .cu_axi10_arqos   (),
  .cu_axi10_arregion(),
  //.cu_axi10_bid     (),
  //.cu_axi10_rid     (),

  .cu_axi11_awready (m_axi_awready[11]),
  .cu_axi11_awvalid (m_axi_awvalid[11]),
  .cu_axi11_awaddr  (m_axi_awaddr [11]),
  .cu_axi11_wready  (m_axi_wready [11]),
  .cu_axi11_wvalid  (m_axi_wvalid [11]),
  .cu_axi11_wdata   (m_axi_wdata  [11]),
  .cu_axi11_wstrb   (m_axi_wstrb  [11]),
  .cu_axi11_wlast   (m_axi_wlast  [11]),
  .cu_axi11_bready  (m_axi_bready [11]),
  .cu_axi11_bvalid  (m_axi_bvalid [11]),
  .cu_axi11_bresp   (m_axi_bresp  [11]),
  .cu_axi11_awburst (m_axi_awburst[11]),
  .cu_axi11_awcache (m_axi_awcache[11]),
  .cu_axi11_awlen   (m_axi_awlen  [11]),
  .cu_axi11_awsize  (m_axi_awsize [11]),
  .cu_axi11_arready (m_axi_arready[11]),
  .cu_axi11_arvalid (m_axi_arvalid[11]),
  .cu_axi11_araddr  (m_axi_araddr [11]),
  .cu_axi11_rready  (m_axi_rready [11]),
  .cu_axi11_rvalid  (m_axi_rvalid [11]),
  .cu_axi11_rdata   (m_axi_rdata  [11]),
  .cu_axi11_rlast   (m_axi_rlast  [11]),
  .cu_axi11_rresp   (m_axi_rresp  [11]),
  .cu_axi11_arburst (m_axi_arburst[11]),
  .cu_axi11_arcache (m_axi_arcache[11]),
  .cu_axi11_arlen   (m_axi_arlen  [11]),
  .cu_axi11_arsize  (m_axi_arsize [11]),
  //.cu_axi11_awid    (),
  .cu_axi11_awprot  (),
  .cu_axi11_awlock  (),
  .cu_axi11_awqos   (),
  .cu_axi11_awregion(),
  //.cu_axi11_arid    (),
  .cu_axi11_arprot  (),
  .cu_axi11_arlock  (),
  .cu_axi11_arqos   (),
  .cu_axi11_arregion(),
  //.cu_axi11_bid     (),
  //.cu_axi11_rid     (),

  .cu_axi12_awready (m_axi_awready[12]),
  .cu_axi12_awvalid (m_axi_awvalid[12]),
  .cu_axi12_awaddr  (m_axi_awaddr [12]),
  .cu_axi12_wready  (m_axi_wready [12]),
  .cu_axi12_wvalid  (m_axi_wvalid [12]),
  .cu_axi12_wdata   (m_axi_wdata  [12]),
  .cu_axi12_wstrb   (m_axi_wstrb  [12]),
  .cu_axi12_wlast   (m_axi_wlast  [12]),
  .cu_axi12_bready  (m_axi_bready [12]),
  .cu_axi12_bvalid  (m_axi_bvalid [12]),
  .cu_axi12_bresp   (m_axi_bresp  [12]),
  .cu_axi12_awburst (m_axi_awburst[12]),
  .cu_axi12_awcache (m_axi_awcache[12]),
  .cu_axi12_awlen   (m_axi_awlen  [12]),
  .cu_axi12_awsize  (m_axi_awsize [12]),
  .cu_axi12_arready (m_axi_arready[12]),
  .cu_axi12_arvalid (m_axi_arvalid[12]),
  .cu_axi12_araddr  (m_axi_araddr [12]),
  .cu_axi12_rready  (m_axi_rready [12]),
  .cu_axi12_rvalid  (m_axi_rvalid [12]),
  .cu_axi12_rdata   (m_axi_rdata  [12]),
  .cu_axi12_rlast   (m_axi_rlast  [12]),
  .cu_axi12_rresp   (m_axi_rresp  [12]),
  .cu_axi12_arburst (m_axi_arburst[12]),
  .cu_axi12_arcache (m_axi_arcache[12]),
  .cu_axi12_arlen   (m_axi_arlen  [12]),
  .cu_axi12_arsize  (m_axi_arsize [12]),
  //.cu_axi12_awid    (),
  .cu_axi12_awprot  (),
  .cu_axi12_awlock  (),
  .cu_axi12_awqos   (),
  .cu_axi12_awregion(),
  //.cu_axi12_arid    (),
  .cu_axi12_arprot  (),
  .cu_axi12_arlock  (),
  .cu_axi12_arqos   (),
  .cu_axi12_arregion(),
  //.cu_axi12_bid     (),
  //.cu_axi12_rid     (),

  .cu_axi13_awready (m_axi_awready[13]),
  .cu_axi13_awvalid (m_axi_awvalid[13]),
  .cu_axi13_awaddr  (m_axi_awaddr [13]),
  .cu_axi13_wready  (m_axi_wready [13]),
  .cu_axi13_wvalid  (m_axi_wvalid [13]),
  .cu_axi13_wdata   (m_axi_wdata  [13]),
  .cu_axi13_wstrb   (m_axi_wstrb  [13]),
  .cu_axi13_wlast   (m_axi_wlast  [13]),
  .cu_axi13_bready  (m_axi_bready [13]),
  .cu_axi13_bvalid  (m_axi_bvalid [13]),
  .cu_axi13_bresp   (m_axi_bresp  [13]),
  .cu_axi13_awburst (m_axi_awburst[13]),
  .cu_axi13_awcache (m_axi_awcache[13]),
  .cu_axi13_awlen   (m_axi_awlen  [13]),
  .cu_axi13_awsize  (m_axi_awsize [13]),
  .cu_axi13_arready (m_axi_arready[13]),
  .cu_axi13_arvalid (m_axi_arvalid[13]),
  .cu_axi13_araddr  (m_axi_araddr [13]),
  .cu_axi13_rready  (m_axi_rready [13]),
  .cu_axi13_rvalid  (m_axi_rvalid [13]),
  .cu_axi13_rdata   (m_axi_rdata  [13]),
  .cu_axi13_rlast   (m_axi_rlast  [13]),
  .cu_axi13_rresp   (m_axi_rresp  [13]),
  .cu_axi13_arburst (m_axi_arburst[13]),
  .cu_axi13_arcache (m_axi_arcache[13]),
  .cu_axi13_arlen   (m_axi_arlen  [13]),
  .cu_axi13_arsize  (m_axi_arsize [13]),
  //.cu_axi13_awid    (),
  .cu_axi13_awprot  (),
  .cu_axi13_awlock  (),
  .cu_axi13_awqos   (),
  .cu_axi13_awregion(),
  //.cu_axi13_arid    (),
  .cu_axi13_arprot  (),
  .cu_axi13_arlock  (),
  .cu_axi13_arqos   (),
  .cu_axi13_arregion(),
  //.cu_axi13_bid     (),
  //.cu_axi13_rid     (),

  .cu_axi14_awready (m_axi_awready[14]),
  .cu_axi14_awvalid (m_axi_awvalid[14]),
  .cu_axi14_awaddr  (m_axi_awaddr [14]),
  .cu_axi14_wready  (m_axi_wready [14]),
  .cu_axi14_wvalid  (m_axi_wvalid [14]),
  .cu_axi14_wdata   (m_axi_wdata  [14]),
  .cu_axi14_wstrb   (m_axi_wstrb  [14]),
  .cu_axi14_wlast   (m_axi_wlast  [14]),
  .cu_axi14_bready  (m_axi_bready [14]),
  .cu_axi14_bvalid  (m_axi_bvalid [14]),
  .cu_axi14_bresp   (m_axi_bresp  [14]),
  .cu_axi14_awburst (m_axi_awburst[14]),
  .cu_axi14_awcache (m_axi_awcache[14]),
  .cu_axi14_awlen   (m_axi_awlen  [14]),
  .cu_axi14_awsize  (m_axi_awsize [14]),
  .cu_axi14_arready (m_axi_arready[14]),
  .cu_axi14_arvalid (m_axi_arvalid[14]),
  .cu_axi14_araddr  (m_axi_araddr [14]),
  .cu_axi14_rready  (m_axi_rready [14]),
  .cu_axi14_rvalid  (m_axi_rvalid [14]),
  .cu_axi14_rdata   (m_axi_rdata  [14]),
  .cu_axi14_rlast   (m_axi_rlast  [14]),
  .cu_axi14_rresp   (m_axi_rresp  [14]),
  .cu_axi14_arburst (m_axi_arburst[14]),
  .cu_axi14_arcache (m_axi_arcache[14]),
  .cu_axi14_arlen   (m_axi_arlen  [14]),
  .cu_axi14_arsize  (m_axi_arsize [14]),
  //.cu_axi14_awid    (),
  .cu_axi14_awprot  (),
  .cu_axi14_awlock  (),
  .cu_axi14_awqos   (),
  .cu_axi14_awregion(),
  //.cu_axi14_arid    (),
  .cu_axi14_arprot  (),
  .cu_axi14_arlock  (),
  .cu_axi14_arqos   (),
  .cu_axi14_arregion(),
  //.cu_axi14_bid     (),
  //.cu_axi14_rid     (),

  .cu_axi15_awready (m_axi_awready[15]),
  .cu_axi15_awvalid (m_axi_awvalid[15]),
  .cu_axi15_awaddr  (m_axi_awaddr [15]),
  .cu_axi15_wready  (m_axi_wready [15]),
  .cu_axi15_wvalid  (m_axi_wvalid [15]),
  .cu_axi15_wdata   (m_axi_wdata  [15]),
  .cu_axi15_wstrb   (m_axi_wstrb  [15]),
  .cu_axi15_wlast   (m_axi_wlast  [15]),
  .cu_axi15_bready  (m_axi_bready [15]),
  .cu_axi15_bvalid  (m_axi_bvalid [15]),
  .cu_axi15_bresp   (m_axi_bresp  [15]),
  .cu_axi15_awburst (m_axi_awburst[15]),
  .cu_axi15_awcache (m_axi_awcache[15]),
  .cu_axi15_awlen   (m_axi_awlen  [15]),
  .cu_axi15_awsize  (m_axi_awsize [15]),
  .cu_axi15_arready (m_axi_arready[15]),
  .cu_axi15_arvalid (m_axi_arvalid[15]),
  .cu_axi15_araddr  (m_axi_araddr [15]),
  .cu_axi15_rready  (m_axi_rready [15]),
  .cu_axi15_rvalid  (m_axi_rvalid [15]),
  .cu_axi15_rdata   (m_axi_rdata  [15]),
  .cu_axi15_rlast   (m_axi_rlast  [15]),
  .cu_axi15_rresp   (m_axi_rresp  [15]),
  .cu_axi15_arburst (m_axi_arburst[15]),
  .cu_axi15_arcache (m_axi_arcache[15]),
  .cu_axi15_arlen   (m_axi_arlen  [15]),
  .cu_axi15_arsize  (m_axi_arsize [15]),
  //.cu_axi15_awid    (),
  .cu_axi15_awprot  (),
  .cu_axi15_awlock  (),
  .cu_axi15_awqos   (),
  .cu_axi15_awregion(),
  //.cu_axi15_arid    (),
  .cu_axi15_arprot  (),
  .cu_axi15_arlock  (),
  .cu_axi15_arqos   (),
  .cu_axi15_arregion()
  //.cu_axi15_bid     (),
  //.cu_axi15_rid     ()
);

`else
bram_init0 bram0 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[0]),
  .s_axi_awvalid(m_axi_awvalid[0]),
  .s_axi_awaddr (m_axi_awaddr [0]),
  .s_axi_wready (m_axi_wready [0]),
  .s_axi_wvalid (m_axi_wvalid [0]),
  .s_axi_wdata  (m_axi_wdata  [0]),
  .s_axi_wstrb  (m_axi_wstrb  [0]),
  .s_axi_wlast  (m_axi_wlast  [0]),
  .s_axi_bready (m_axi_bready [0]),
  .s_axi_bvalid (m_axi_bvalid [0]),
  .s_axi_bresp  (m_axi_bresp  [0]),
  .s_axi_awlen  (m_axi_awlen  [0]),
  .s_axi_awsize (m_axi_awsize [0]),
  .s_axi_awburst(m_axi_awburst[0]),
  .s_axi_arready(m_axi_arready[0]),
  .s_axi_arvalid(m_axi_arvalid[0]),
  .s_axi_araddr (m_axi_araddr [0]),
  .s_axi_rready (m_axi_rready [0]),
  .s_axi_rvalid (m_axi_rvalid [0]),
  .s_axi_rdata  (m_axi_rdata  [0]),
  .s_axi_rlast  (m_axi_rlast  [0]),
  .s_axi_rresp  (m_axi_rresp  [0]),
  .s_axi_arlen  (m_axi_arlen  [0]),
  .s_axi_arsize (m_axi_arsize [0]),
  .s_axi_arburst(m_axi_arburst[0]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init1 bram1 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[1]),
  .s_axi_awvalid(m_axi_awvalid[1]),
  .s_axi_awaddr (m_axi_awaddr [1]),
  .s_axi_wready (m_axi_wready [1]),
  .s_axi_wvalid (m_axi_wvalid [1]),
  .s_axi_wdata  (m_axi_wdata  [1]),
  .s_axi_wstrb  (m_axi_wstrb  [1]),
  .s_axi_wlast  (m_axi_wlast  [1]),
  .s_axi_bready (m_axi_bready [1]),
  .s_axi_bvalid (m_axi_bvalid [1]),
  .s_axi_bresp  (m_axi_bresp  [1]),
  .s_axi_awlen  (m_axi_awlen  [1]),
  .s_axi_awsize (m_axi_awsize [1]),
  .s_axi_awburst(m_axi_awburst[1]),
  .s_axi_arready(m_axi_arready[1]),
  .s_axi_arvalid(m_axi_arvalid[1]),
  .s_axi_araddr (m_axi_araddr [1]),
  .s_axi_rready (m_axi_rready [1]),
  .s_axi_rvalid (m_axi_rvalid [1]),
  .s_axi_rdata  (m_axi_rdata  [1]),
  .s_axi_rlast  (m_axi_rlast  [1]),
  .s_axi_rresp  (m_axi_rresp  [1]),
  .s_axi_arlen  (m_axi_arlen  [1]),
  .s_axi_arsize (m_axi_arsize [1]),
  .s_axi_arburst(m_axi_arburst[1]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init2 bram2 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[2]),
  .s_axi_awvalid(m_axi_awvalid[2]),
  .s_axi_awaddr (m_axi_awaddr [2]),
  .s_axi_wready (m_axi_wready [2]),
  .s_axi_wvalid (m_axi_wvalid [2]),
  .s_axi_wdata  (m_axi_wdata  [2]),
  .s_axi_wstrb  (m_axi_wstrb  [2]),
  .s_axi_wlast  (m_axi_wlast  [2]),
  .s_axi_bready (m_axi_bready [2]),
  .s_axi_bvalid (m_axi_bvalid [2]),
  .s_axi_bresp  (m_axi_bresp  [2]),
  .s_axi_awlen  (m_axi_awlen  [2]),
  .s_axi_awsize (m_axi_awsize [2]),
  .s_axi_awburst(m_axi_awburst[2]),
  .s_axi_arready(m_axi_arready[2]),
  .s_axi_arvalid(m_axi_arvalid[2]),
  .s_axi_araddr (m_axi_araddr [2]),
  .s_axi_rready (m_axi_rready [2]),
  .s_axi_rvalid (m_axi_rvalid [2]),
  .s_axi_rdata  (m_axi_rdata  [2]),
  .s_axi_rlast  (m_axi_rlast  [2]),
  .s_axi_rresp  (m_axi_rresp  [2]),
  .s_axi_arlen  (m_axi_arlen  [2]),
  .s_axi_arsize (m_axi_arsize [2]),
  .s_axi_arburst(m_axi_arburst[2]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init3 bram3 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[3]),
  .s_axi_awvalid(m_axi_awvalid[3]),
  .s_axi_awaddr (m_axi_awaddr [3]),
  .s_axi_wready (m_axi_wready [3]),
  .s_axi_wvalid (m_axi_wvalid [3]),
  .s_axi_wdata  (m_axi_wdata  [3]),
  .s_axi_wstrb  (m_axi_wstrb  [3]),
  .s_axi_wlast  (m_axi_wlast  [3]),
  .s_axi_bready (m_axi_bready [3]),
  .s_axi_bvalid (m_axi_bvalid [3]),
  .s_axi_bresp  (m_axi_bresp  [3]),
  .s_axi_awlen  (m_axi_awlen  [3]),
  .s_axi_awsize (m_axi_awsize [3]),
  .s_axi_awburst(m_axi_awburst[3]),
  .s_axi_arready(m_axi_arready[3]),
  .s_axi_arvalid(m_axi_arvalid[3]),
  .s_axi_araddr (m_axi_araddr [3]),
  .s_axi_rready (m_axi_rready [3]),
  .s_axi_rvalid (m_axi_rvalid [3]),
  .s_axi_rdata  (m_axi_rdata  [3]),
  .s_axi_rlast  (m_axi_rlast  [3]),
  .s_axi_rresp  (m_axi_rresp  [3]),
  .s_axi_arlen  (m_axi_arlen  [3]),
  .s_axi_arsize (m_axi_arsize [3]),
  .s_axi_arburst(m_axi_arburst[3]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init4 bram4 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[4]),
  .s_axi_awvalid(m_axi_awvalid[4]),
  .s_axi_awaddr (m_axi_awaddr [4]),
  .s_axi_wready (m_axi_wready [4]),
  .s_axi_wvalid (m_axi_wvalid [4]),
  .s_axi_wdata  (m_axi_wdata  [4]),
  .s_axi_wstrb  (m_axi_wstrb  [4]),
  .s_axi_wlast  (m_axi_wlast  [4]),
  .s_axi_bready (m_axi_bready [4]),
  .s_axi_bvalid (m_axi_bvalid [4]),
  .s_axi_bresp  (m_axi_bresp  [4]),
  .s_axi_awlen  (m_axi_awlen  [4]),
  .s_axi_awsize (m_axi_awsize [4]),
  .s_axi_awburst(m_axi_awburst[4]),
  .s_axi_arready(m_axi_arready[4]),
  .s_axi_arvalid(m_axi_arvalid[4]),
  .s_axi_araddr (m_axi_araddr [4]),
  .s_axi_rready (m_axi_rready [4]),
  .s_axi_rvalid (m_axi_rvalid [4]),
  .s_axi_rdata  (m_axi_rdata  [4]),
  .s_axi_rlast  (m_axi_rlast  [4]),
  .s_axi_rresp  (m_axi_rresp  [4]),
  .s_axi_arlen  (m_axi_arlen  [4]),
  .s_axi_arsize (m_axi_arsize [4]),
  .s_axi_arburst(m_axi_arburst[4]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init5 bram5 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[5]),
  .s_axi_awvalid(m_axi_awvalid[5]),
  .s_axi_awaddr (m_axi_awaddr [5]),
  .s_axi_wready (m_axi_wready [5]),
  .s_axi_wvalid (m_axi_wvalid [5]),
  .s_axi_wdata  (m_axi_wdata  [5]),
  .s_axi_wstrb  (m_axi_wstrb  [5]),
  .s_axi_wlast  (m_axi_wlast  [5]),
  .s_axi_bready (m_axi_bready [5]),
  .s_axi_bvalid (m_axi_bvalid [5]),
  .s_axi_bresp  (m_axi_bresp  [5]),
  .s_axi_awlen  (m_axi_awlen  [5]),
  .s_axi_awsize (m_axi_awsize [5]),
  .s_axi_awburst(m_axi_awburst[5]),
  .s_axi_arready(m_axi_arready[5]),
  .s_axi_arvalid(m_axi_arvalid[5]),
  .s_axi_araddr (m_axi_araddr [5]),
  .s_axi_rready (m_axi_rready [5]),
  .s_axi_rvalid (m_axi_rvalid [5]),
  .s_axi_rdata  (m_axi_rdata  [5]),
  .s_axi_rlast  (m_axi_rlast  [5]),
  .s_axi_rresp  (m_axi_rresp  [5]),
  .s_axi_arlen  (m_axi_arlen  [5]),
  .s_axi_arsize (m_axi_arsize [5]),
  .s_axi_arburst(m_axi_arburst[5]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init6 bram6 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[6]),
  .s_axi_awvalid(m_axi_awvalid[6]),
  .s_axi_awaddr (m_axi_awaddr [6]),
  .s_axi_wready (m_axi_wready [6]),
  .s_axi_wvalid (m_axi_wvalid [6]),
  .s_axi_wdata  (m_axi_wdata  [6]),
  .s_axi_wstrb  (m_axi_wstrb  [6]),
  .s_axi_wlast  (m_axi_wlast  [6]),
  .s_axi_bready (m_axi_bready [6]),
  .s_axi_bvalid (m_axi_bvalid [6]),
  .s_axi_bresp  (m_axi_bresp  [6]),
  .s_axi_awlen  (m_axi_awlen  [6]),
  .s_axi_awsize (m_axi_awsize [6]),
  .s_axi_awburst(m_axi_awburst[6]),
  .s_axi_arready(m_axi_arready[6]),
  .s_axi_arvalid(m_axi_arvalid[6]),
  .s_axi_araddr (m_axi_araddr [6]),
  .s_axi_rready (m_axi_rready [6]),
  .s_axi_rvalid (m_axi_rvalid [6]),
  .s_axi_rdata  (m_axi_rdata  [6]),
  .s_axi_rlast  (m_axi_rlast  [6]),
  .s_axi_rresp  (m_axi_rresp  [6]),
  .s_axi_arlen  (m_axi_arlen  [6]),
  .s_axi_arsize (m_axi_arsize [6]),
  .s_axi_arburst(m_axi_arburst[6]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init7 bram7 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[7]),
  .s_axi_awvalid(m_axi_awvalid[7]),
  .s_axi_awaddr (m_axi_awaddr [7]),
  .s_axi_wready (m_axi_wready [7]),
  .s_axi_wvalid (m_axi_wvalid [7]),
  .s_axi_wdata  (m_axi_wdata  [7]),
  .s_axi_wstrb  (m_axi_wstrb  [7]),
  .s_axi_wlast  (m_axi_wlast  [7]),
  .s_axi_bready (m_axi_bready [7]),
  .s_axi_bvalid (m_axi_bvalid [7]),
  .s_axi_bresp  (m_axi_bresp  [7]),
  .s_axi_awlen  (m_axi_awlen  [7]),
  .s_axi_awsize (m_axi_awsize [7]),
  .s_axi_awburst(m_axi_awburst[7]),
  .s_axi_arready(m_axi_arready[7]),
  .s_axi_arvalid(m_axi_arvalid[7]),
  .s_axi_araddr (m_axi_araddr [7]),
  .s_axi_rready (m_axi_rready [7]),
  .s_axi_rvalid (m_axi_rvalid [7]),
  .s_axi_rdata  (m_axi_rdata  [7]),
  .s_axi_rlast  (m_axi_rlast  [7]),
  .s_axi_rresp  (m_axi_rresp  [7]),
  .s_axi_arlen  (m_axi_arlen  [7]),
  .s_axi_arsize (m_axi_arsize [7]),
  .s_axi_arburst(m_axi_arburst[7]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init8 bram8 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[8]),
  .s_axi_awvalid(m_axi_awvalid[8]),
  .s_axi_awaddr (m_axi_awaddr [8]),
  .s_axi_wready (m_axi_wready [8]),
  .s_axi_wvalid (m_axi_wvalid [8]),
  .s_axi_wdata  (m_axi_wdata  [8]),
  .s_axi_wstrb  (m_axi_wstrb  [8]),
  .s_axi_wlast  (m_axi_wlast  [8]),
  .s_axi_bready (m_axi_bready [8]),
  .s_axi_bvalid (m_axi_bvalid [8]),
  .s_axi_bresp  (m_axi_bresp  [8]),
  .s_axi_awlen  (m_axi_awlen  [8]),
  .s_axi_awsize (m_axi_awsize [8]),
  .s_axi_awburst(m_axi_awburst[8]),
  .s_axi_arready(m_axi_arready[8]),
  .s_axi_arvalid(m_axi_arvalid[8]),
  .s_axi_araddr (m_axi_araddr [8]),
  .s_axi_rready (m_axi_rready [8]),
  .s_axi_rvalid (m_axi_rvalid [8]),
  .s_axi_rdata  (m_axi_rdata  [8]),
  .s_axi_rlast  (m_axi_rlast  [8]),
  .s_axi_rresp  (m_axi_rresp  [8]),
  .s_axi_arlen  (m_axi_arlen  [8]),
  .s_axi_arsize (m_axi_arsize [8]),
  .s_axi_arburst(m_axi_arburst[8]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init9 bram9 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[9]),
  .s_axi_awvalid(m_axi_awvalid[9]),
  .s_axi_awaddr (m_axi_awaddr [9]),
  .s_axi_wready (m_axi_wready [9]),
  .s_axi_wvalid (m_axi_wvalid [9]),
  .s_axi_wdata  (m_axi_wdata  [9]),
  .s_axi_wstrb  (m_axi_wstrb  [9]),
  .s_axi_wlast  (m_axi_wlast  [9]),
  .s_axi_bready (m_axi_bready [9]),
  .s_axi_bvalid (m_axi_bvalid [9]),
  .s_axi_bresp  (m_axi_bresp  [9]),
  .s_axi_awlen  (m_axi_awlen  [9]),
  .s_axi_awsize (m_axi_awsize [9]),
  .s_axi_awburst(m_axi_awburst[9]),
  .s_axi_arready(m_axi_arready[9]),
  .s_axi_arvalid(m_axi_arvalid[9]),
  .s_axi_araddr (m_axi_araddr [9]),
  .s_axi_rready (m_axi_rready [9]),
  .s_axi_rvalid (m_axi_rvalid [9]),
  .s_axi_rdata  (m_axi_rdata  [9]),
  .s_axi_rlast  (m_axi_rlast  [9]),
  .s_axi_rresp  (m_axi_rresp  [9]),
  .s_axi_arlen  (m_axi_arlen  [9]),
  .s_axi_arsize (m_axi_arsize [9]),
  .s_axi_arburst(m_axi_arburst[9]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init10 bram10 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[10]),
  .s_axi_awvalid(m_axi_awvalid[10]),
  .s_axi_awaddr (m_axi_awaddr [10]),
  .s_axi_wready (m_axi_wready [10]),
  .s_axi_wvalid (m_axi_wvalid [10]),
  .s_axi_wdata  (m_axi_wdata  [10]),
  .s_axi_wstrb  (m_axi_wstrb  [10]),
  .s_axi_wlast  (m_axi_wlast  [10]),
  .s_axi_bready (m_axi_bready [10]),
  .s_axi_bvalid (m_axi_bvalid [10]),
  .s_axi_bresp  (m_axi_bresp  [10]),
  .s_axi_awlen  (m_axi_awlen  [10]),
  .s_axi_awsize (m_axi_awsize [10]),
  .s_axi_awburst(m_axi_awburst[10]),
  .s_axi_arready(m_axi_arready[10]),
  .s_axi_arvalid(m_axi_arvalid[10]),
  .s_axi_araddr (m_axi_araddr [10]),
  .s_axi_rready (m_axi_rready [10]),
  .s_axi_rvalid (m_axi_rvalid [10]),
  .s_axi_rdata  (m_axi_rdata  [10]),
  .s_axi_rlast  (m_axi_rlast  [10]),
  .s_axi_rresp  (m_axi_rresp  [10]),
  .s_axi_arlen  (m_axi_arlen  [10]),
  .s_axi_arsize (m_axi_arsize [10]),
  .s_axi_arburst(m_axi_arburst[10]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init11 bram11 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[11]),
  .s_axi_awvalid(m_axi_awvalid[11]),
  .s_axi_awaddr (m_axi_awaddr [11]),
  .s_axi_wready (m_axi_wready [11]),
  .s_axi_wvalid (m_axi_wvalid [11]),
  .s_axi_wdata  (m_axi_wdata  [11]),
  .s_axi_wstrb  (m_axi_wstrb  [11]),
  .s_axi_wlast  (m_axi_wlast  [11]),
  .s_axi_bready (m_axi_bready [11]),
  .s_axi_bvalid (m_axi_bvalid [11]),
  .s_axi_bresp  (m_axi_bresp  [11]),
  .s_axi_awlen  (m_axi_awlen  [11]),
  .s_axi_awsize (m_axi_awsize [11]),
  .s_axi_awburst(m_axi_awburst[11]),
  .s_axi_arready(m_axi_arready[11]),
  .s_axi_arvalid(m_axi_arvalid[11]),
  .s_axi_araddr (m_axi_araddr [11]),
  .s_axi_rready (m_axi_rready [11]),
  .s_axi_rvalid (m_axi_rvalid [11]),
  .s_axi_rdata  (m_axi_rdata  [11]),
  .s_axi_rlast  (m_axi_rlast  [11]),
  .s_axi_rresp  (m_axi_rresp  [11]),
  .s_axi_arlen  (m_axi_arlen  [11]),
  .s_axi_arsize (m_axi_arsize [11]),
  .s_axi_arburst(m_axi_arburst[11]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init12 bram12 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[12]),
  .s_axi_awvalid(m_axi_awvalid[12]),
  .s_axi_awaddr (m_axi_awaddr [12]),
  .s_axi_wready (m_axi_wready [12]),
  .s_axi_wvalid (m_axi_wvalid [12]),
  .s_axi_wdata  (m_axi_wdata  [12]),
  .s_axi_wstrb  (m_axi_wstrb  [12]),
  .s_axi_wlast  (m_axi_wlast  [12]),
  .s_axi_bready (m_axi_bready [12]),
  .s_axi_bvalid (m_axi_bvalid [12]),
  .s_axi_bresp  (m_axi_bresp  [12]),
  .s_axi_awlen  (m_axi_awlen  [12]),
  .s_axi_awsize (m_axi_awsize [12]),
  .s_axi_awburst(m_axi_awburst[12]),
  .s_axi_arready(m_axi_arready[12]),
  .s_axi_arvalid(m_axi_arvalid[12]),
  .s_axi_araddr (m_axi_araddr [12]),
  .s_axi_rready (m_axi_rready [12]),
  .s_axi_rvalid (m_axi_rvalid [12]),
  .s_axi_rdata  (m_axi_rdata  [12]),
  .s_axi_rlast  (m_axi_rlast  [12]),
  .s_axi_rresp  (m_axi_rresp  [12]),
  .s_axi_arlen  (m_axi_arlen  [12]),
  .s_axi_arsize (m_axi_arsize [12]),
  .s_axi_arburst(m_axi_arburst[12]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init13 bram13 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[13]),
  .s_axi_awvalid(m_axi_awvalid[13]),
  .s_axi_awaddr (m_axi_awaddr [13]),
  .s_axi_wready (m_axi_wready [13]),
  .s_axi_wvalid (m_axi_wvalid [13]),
  .s_axi_wdata  (m_axi_wdata  [13]),
  .s_axi_wstrb  (m_axi_wstrb  [13]),
  .s_axi_wlast  (m_axi_wlast  [13]),
  .s_axi_bready (m_axi_bready [13]),
  .s_axi_bvalid (m_axi_bvalid [13]),
  .s_axi_bresp  (m_axi_bresp  [13]),
  .s_axi_awlen  (m_axi_awlen  [13]),
  .s_axi_awsize (m_axi_awsize [13]),
  .s_axi_awburst(m_axi_awburst[13]),
  .s_axi_arready(m_axi_arready[13]),
  .s_axi_arvalid(m_axi_arvalid[13]),
  .s_axi_araddr (m_axi_araddr [13]),
  .s_axi_rready (m_axi_rready [13]),
  .s_axi_rvalid (m_axi_rvalid [13]),
  .s_axi_rdata  (m_axi_rdata  [13]),
  .s_axi_rlast  (m_axi_rlast  [13]),
  .s_axi_rresp  (m_axi_rresp  [13]),
  .s_axi_arlen  (m_axi_arlen  [13]),
  .s_axi_arsize (m_axi_arsize [13]),
  .s_axi_arburst(m_axi_arburst[13]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init14 bram14 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[14]),
  .s_axi_awvalid(m_axi_awvalid[14]),
  .s_axi_awaddr (m_axi_awaddr [14]),
  .s_axi_wready (m_axi_wready [14]),
  .s_axi_wvalid (m_axi_wvalid [14]),
  .s_axi_wdata  (m_axi_wdata  [14]),
  .s_axi_wstrb  (m_axi_wstrb  [14]),
  .s_axi_wlast  (m_axi_wlast  [14]),
  .s_axi_bready (m_axi_bready [14]),
  .s_axi_bvalid (m_axi_bvalid [14]),
  .s_axi_bresp  (m_axi_bresp  [14]),
  .s_axi_awlen  (m_axi_awlen  [14]),
  .s_axi_awsize (m_axi_awsize [14]),
  .s_axi_awburst(m_axi_awburst[14]),
  .s_axi_arready(m_axi_arready[14]),
  .s_axi_arvalid(m_axi_arvalid[14]),
  .s_axi_araddr (m_axi_araddr [14]),
  .s_axi_rready (m_axi_rready [14]),
  .s_axi_rvalid (m_axi_rvalid [14]),
  .s_axi_rdata  (m_axi_rdata  [14]),
  .s_axi_rlast  (m_axi_rlast  [14]),
  .s_axi_rresp  (m_axi_rresp  [14]),
  .s_axi_arlen  (m_axi_arlen  [14]),
  .s_axi_arsize (m_axi_arsize [14]),
  .s_axi_arburst(m_axi_arburst[14]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init15 bram15 (
  .s_aclk       (sclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(m_axi_awready[15]),
  .s_axi_awvalid(m_axi_awvalid[15]),
  .s_axi_awaddr (m_axi_awaddr [15]),
  .s_axi_wready (m_axi_wready [15]),
  .s_axi_wvalid (m_axi_wvalid [15]),
  .s_axi_wdata  (m_axi_wdata  [15]),
  .s_axi_wstrb  (m_axi_wstrb  [15]),
  .s_axi_wlast  (m_axi_wlast  [15]),
  .s_axi_bready (m_axi_bready [15]),
  .s_axi_bvalid (m_axi_bvalid [15]),
  .s_axi_bresp  (m_axi_bresp  [15]),
  .s_axi_awlen  (m_axi_awlen  [15]),
  .s_axi_awsize (m_axi_awsize [15]),
  .s_axi_awburst(m_axi_awburst[15]),
  .s_axi_arready(m_axi_arready[15]),
  .s_axi_arvalid(m_axi_arvalid[15]),
  .s_axi_araddr (m_axi_araddr [15]),
  .s_axi_rready (m_axi_rready [15]),
  .s_axi_rvalid (m_axi_rvalid [15]),
  .s_axi_rdata  (m_axi_rdata  [15]),
  .s_axi_rlast  (m_axi_rlast  [15]),
  .s_axi_rresp  (m_axi_rresp  [15]),
  .s_axi_arlen  (m_axi_arlen  [15]),
  .s_axi_arsize (m_axi_arsize [15]),
  .s_axi_arburst(m_axi_arburst[15]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);
`endif

wire [NUM_GROUP-1:0] launch;
wire [NUM_GROUP-1:0] start_load;
inte #(
  .NUM_GROUP(NUM_GROUP)
) inte_i (
  .sclk          (sclk),
  .xdma_rstn     (xdma_rstn),
  .gpio          (gpio),
  .start_load    (start_load),
  .rst_n         (rst_n),
  .launch        (launch),
  .start_load_all(start_load_all)
);

/**************************** 数据加载 ****************************/
wire   [NUM_GROUP-1:0] start_turn;
wire   [NUM_GROUP-1:0] done_upload;
wire   [NUM_GROUP-1:0] upload;
wire  [SIZE_GROUP-1:0] wea_load   [NUM_GROUP-1:0];
wire [AWIDTH_BRAM-1:0] addra_load [NUM_GROUP-1:0];
wire [AWIDTH_BRAM-1:0] addrb_load [NUM_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] dout_load  [NUM_GROUP-1:0][SIZE_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] din_load   [NUM_GROUP-1:0][SIZE_GROUP-1:0];
assign upload = start_load; 
generate for (genvar m=0; m<NUM_GROUP; m=m+1) begin
  load #(
    .ID_GROUP   (m),
    .LENGTH     (LENGTH),
    .SIZE_LOOP  (SIZE_LOOP),
    .SIZE_GROUP (SIZE_GROUP),
    .AWIDTH_HBM (AWIDTH_HBM),
    .DWIDTH_HBM (DWIDTH_HBM),
    .DWIDTH_BRAM(DWIDTH_BRAM),
    .AWIDTH_BRAM(AWIDTH_BRAM)
  ) load_i (
    .sclk        (sclk),
    .rst_n       (rst_n),
    .launch      (launch[m]),
    .wea_load    (wea_load[m]),
    .addra_load  (addra_load[m]),
    .addrb_load  (addrb_load[m]),
    .start_load  (start_load[m]),
    .upload      (upload[m]),
    .done_upload (done_upload[m]),

    .dout_load0  (dout_load[m][0]),
    .dout_load1  (dout_load[m][1]),
    .dout_load2  (dout_load[m][2]),
    .dout_load3  (dout_load[m][3]),
    .dout_load4  (dout_load[m][4]),
    .dout_load5  (dout_load[m][5]),
    .dout_load6  (dout_load[m][6]),
    .dout_load7  (dout_load[m][7]),

    .din_load0  (din_load[m][0]),
    .din_load1  (din_load[m][1]),
    .din_load2  (din_load[m][2]),
    .din_load3  (din_load[m][3]),
    .din_load4  (din_load[m][4]),
    .din_load5  (din_load[m][5]),
    .din_load6  (din_load[m][6]),
    .din_load7  (din_load[m][7]),

    .axi_awready(m_axi_awready[m]),
    .axi_awvalid(m_axi_awvalid[m]),
    .axi_awaddr (m_axi_awaddr [m]),
    .axi_awburst(m_axi_awburst[m]),
    .axi_awlen  (m_axi_awlen  [m]),
    .axi_awcache(m_axi_awcache[m]),
    .axi_awsize (m_axi_awsize [m]),
    .axi_wready (m_axi_wready [m]),
    .axi_wvalid (m_axi_wvalid [m]),
    .axi_wdata  (m_axi_wdata  [m]),
    .axi_wstrb  (m_axi_wstrb  [m]),
    .axi_wlast  (m_axi_wlast  [m]),
    .axi_bready (m_axi_bready [m]),
    .axi_bvalid (m_axi_bvalid [m]),
    .axi_bresp  (m_axi_bresp  [m]),
    .axi_arready(m_axi_arready[m]),
    .axi_arvalid(m_axi_arvalid[m]),
    .axi_araddr (m_axi_araddr [m]),
    .axi_arburst(m_axi_arburst[m]),
    .axi_arlen  (m_axi_arlen  [m]),
    .axi_arcache(m_axi_arcache[m]),
    .axi_arsize (m_axi_arsize [m]),
    .axi_rready (m_axi_rready [m]),
    .axi_rvalid (m_axi_rvalid [m]),
    .axi_rdata  (m_axi_rdata  [m]),
    .axi_rlast  (m_axi_rlast  [m]),
    .axi_rresp  (m_axi_rresp  [m])
  );
end
endgenerate

/**************************** 数据缓存 ****************************/
wire   [NUM_GROUP-1:0] web_sw ;
wire [AWIDTH_BRAM-1:0] addrb_sw  [NUM_GROUP-1:0];
wire [AWIDTH_BRAM-1:0] addrb_fft [NUM_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] din_fft   [NUM_GROUP-1:0][SIZE_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] dout_sw   [NUM_GROUP-1:0][SIZE_GROUP-1:0];
generate for (genvar m=0; m<NUM_GROUP; m=m+1) begin
mem #(
  .ID_GROUP   (m),
  .LENGTH     (LENGTH),
  .SIZE_LOOP  (SIZE_LOOP),
  .SIZE_GROUP (SIZE_GROUP),
  .DWIDTH_BRAM(DWIDTH_BRAM),
  .AWIDTH_BRAM(AWIDTH_BRAM)
) mem_i (
  .sclk   (sclk),
  .rst_n  (rst_n),
  .flag0  (0),
  .flag1  (0),

  .wea    (wea_load[m]),
  .addra  (addra_load[m]),
  .dina0  (dout_load[m][0]),
  .dina1  (dout_load[m][1]),
  .dina2  (dout_load[m][2]),
  .dina3  (dout_load[m][3]),
  .dina4  (dout_load[m][4]),
  .dina5  (dout_load[m][5]),
  .dina6  (dout_load[m][6]),
  .dina7  (dout_load[m][7]),

  .web    (web_sw[m]),
  .addrb  (addrb_sw[m]),
  .dinb0  (dout_sw[m][0]),
  .dinb1  (dout_sw[m][1]),
  .dinb2  (dout_sw[m][2]),
  .dinb3  (dout_sw[m][3]),
  .dinb4  (dout_sw[m][4]),
  .dinb5  (dout_sw[m][5]),
  .dinb6  (dout_sw[m][6]),
  .dinb7  (dout_sw[m][7]),

  .addrc  (addrb_load[m]),
  .douta0 (din_load[m][0]),
  .douta1 (din_load[m][1]),
  .douta2 (din_load[m][2]),
  .douta3 (din_load[m][3]),
  .douta4 (din_load[m][4]),
  .douta5 (din_load[m][5]),
  .douta6 (din_load[m][6]),
  .douta7 (din_load[m][7]),

  .addrd  (addrb_fft[m]),
  .doutb0 (din_fft[m][0]),
  .doutb1 (din_fft[m][1]),
  .doutb2 (din_fft[m][2]),
  .doutb3 (din_fft[m][3]),
  .doutb4 (din_fft[m][4]),
  .doutb5 (din_fft[m][5]),
  .doutb6 (din_fft[m][6]),
  .doutb7 (din_fft[m][7])
);
end
endgenerate

/**************************** 数据监控 ****************************/
ila ila_i (
  .clk(sclk),
  .probe0 (m_axi_awready[0]),
  .probe1 (m_axi_awvalid[0]),
  .probe2 (m_axi_awaddr [0]),
  .probe3 (m_axi_wready [0]),
  .probe4 (m_axi_wvalid [0]),
  .probe5 (m_axi_wdata  [0]),
  .probe6 (m_axi_wstrb  [0]),
  .probe7 (m_axi_wlast  [0]),
  .probe8 (m_axi_arready[0]),
  .probe9 (m_axi_arvalid[0]),
  .probe10(m_axi_araddr [0]),
  .probe11(m_axi_rready [0]),
  .probe12(m_axi_rvalid [0]),
  .probe13(m_axi_rdata  [0]),
  .probe14(m_axi_rlast  [0]),
  .probe15(m_axi_awready[15]),
  .probe16(m_axi_awvalid[15]),
  .probe17(m_axi_awaddr [15]),
  .probe18(m_axi_wready [15]),
  .probe19(m_axi_wvalid [15]),
  .probe20(m_axi_wdata  [15]),
  .probe21(m_axi_wstrb  [15]),
  .probe22(m_axi_wlast  [15]),
  .probe23(m_axi_arready[15]),
  .probe24(m_axi_arvalid[15]),
  .probe25(m_axi_araddr [15]),
  .probe26(m_axi_rready [15]),
  .probe27(m_axi_rvalid [15]),
  .probe28(m_axi_rdata  [15]),
  .probe29(m_axi_rlast  [15]),
  .probe30(launch           )
);

endmodule