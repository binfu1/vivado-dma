`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NyUsoNEOp4jN8y7wOwKG+OLRKfYfA5+orGMeKd7sK0Mz8f6rkD8Cd4ee5gtDF5WWj3Bbyj/fN7pD
kOIbJEOt9yicq3th7leCwF1FYui+HkOHrAJn82fBKmgsUxAS6zLI2r65N7awfSOXOdUzS9S4iv0j
VnAgQzvmk50i5eOArjtLNGUxiRN5xjmEjNuZ2A/uRVxBM2bSRZvSipyC8vPOCOQd95FFIFg7Oj1D
G2udGUZI+r12yu2ICnkDpIvVrzM1icds5ynCNl6hkJhFiBBwWHnh7btPNA26jAiGAtlY3LdMzMu+
3yfWfZMr8QXEbLyAW/aFBJ4okE+9m7+eqyeSHA==
`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cckiFnXuCWvElG/8IVGT6Uhku1/SgNaWtMSigVERkVYUUbn+DTffLdBCEmtJhkJmZB73lwzNFdaq
7Tl6CUBOU/k3Gus4DzctATBZEYYP5UpDI+gTPvEwNLcR+SyK+rzbgcnzUTb1uiqPKD8/S4a49PEr
R4yJ4w19Z7JneOzXVfr4xIxHyR7C5IMRez94VSWzTanP2ohrOiqdDTkUUA58LUU2dOABnEjEegpv
d7b9FQIU1LeV5Gz6a+TZ95JNQvjfgL2UDWzCKiwHi0X2UbFmSMLbQFAwLQQ4d7BfH3N+N7lmL0FU
CRVrUmNiVJyCZaNGNWP1qAtHyU/3XRxsWmZzLg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
RojZU0NT3tJcOK6vvTGSS/bpgAe+P3EP8USJfiF7t8XLeIcTsNnkba80WrhB867eE/K5TGEFbQed
g0EnBglD2Q==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mfjGCX7fcqP5dTxLxc8xSDcjkpu89+26N8NsThgZL9iWZn7Z3Ygf0KYPmRXzyIWkvtulW3Q+tp1C
Hj+hPyfzZeeyJu/v2BwmBv5oOmJK2/DTnlJA/a+86nu2DslE5CpDoVNB5ASE0/gh94akQcDt4wQe
ORYPCw0L6mDTjlE2vGE5/q6lPSjhtEa/f6M2ud+Y0n6xP5ZJgoFazaw+YCPKhpm8ho8wLZU+ADEW
4nxXH/wfBGjJZQdFiSo6cUySCV3h1faor6fAE5cVxi9ZktW35LmZRts/qJk57z5T0ip2sAtKaIQ+
yOHv9LvZFXZ3MjdiwUM1J7PXB1U5bGIqCKtE1Q==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Oc48AMFGwNE4bxAIFLTq/LsNnFj3/Sha26BoBLJAhsSzsT7xKrHVkCIEMRRp6sUDmyKBthEhUeAZ
u3XRi8E5wqLH6Z6xJ2dYDKkcMEhbjCAMCyGAOnUFWWE3tR4MI6bncFKYLeKwFzjq8wjBlzyvFCNz
3ZfZbzdO1SULnOInCwE=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BFF3tXKXQxNkcfVkkYL6Huk49khrP4/X59P/vVmv5/+M+sTNqmxVEqn+YFlBUzhV9ZKgZD8NCpEj
/XbLGO7gXXDEcaGDsjOjLP7Uj4/AVfQ8dcUw71A19YPFkGzQk3fpS/KvDXVNxEDXXw17tETTCEVf
PnZWFpdpivZWNmYFcIVi+avEPOzRky4KbzBdt6bwziA/TvSa1nSG+U2kDIbhErGyAQUeGfRnRy9X
XNc3hCfvmtcq9q6AqOr7I8fpoUiK7D5ShILguvb7yiZPCUOVrconJGo6UBzIQGktQLATvHqifgVq
globS8t/iEGH9i8hBWKxlPEu2tMYeBypZuGYEA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lEmc+h5qPNSuLjd69zuJzgsK6kqBZxjOCma4OF901m9pDPMrMXhBqg567djgIpEnYZG7Ir2cEW1K
h+JMx5YS2JiI+X4AnbXsTy7cPf3EPLQoQJiYd4z0EVpssmaESSwBpcJHe6xWuZ3jh8a6BZynP80G
7xcTZn/poN7geM4Y4QldbmFR73YKjsOv5rJLj3U3URN2211SSe78WpHvGzx01HIRTgVITvOTGgDI
Mozb5NN+u1dtQIsP97+RHLGkYhA7KcjJXDc7sPcjBUR15RR175W0PDtAwLfeyxW1oEKnSd7AURrD
u5kPjIet80JNcjBGMh3PHlnWBy7drNj84pUV7g==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
g/rneQ4eAHoU68Py3fPvHQVFMAzXaNQOA8DP9q3N6az6xvq/Et5Q3d1n7vmq4cFmTg5eMBPQBnLq
EyfE6TkZYtldzmlWTP641bnhzvrT0SMnfmfJv+9xhGr19Vufp+fIY9+7DZ3lmfuuJ7Ru1kYrgelm
j37qKvBGlOGqyl+vW9s=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GVSlRhl+0id9zKmLY/wvDnOK+m1jWKwawbu6WXASN51dQB904Klo7OvRtTsa9nnAENxUiE8w7OwC
K2GmuKgUKEfVFD/L4TvqPQBByJ43VtRwEIcavzB6v4Wxrbr/ZIxSbkeLDegWAoEwRd5lzUYfK6FE
cC8F6yFhRlnBxPKv8V0gtw/0ulxL7BbxUEwvVARwMXDcHe2qX5yjMdgaZe6xnSV9Ma9W/GO/EAD4
VM8Evr4nMWFueWgv5U7oa07HNa104V2PlB1IDsQiysdkIuNIIRqc2EGkGEAs2x/4pL/mXpMBIbZR
F6Oy6w3e9pFywHsyrt3ZAV01yP6AH3Eb27gsFg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
yuZr0X/f7JxatSvKrNTFABRdsGtu8o7MUgVf1FC7CT++z3U8dkzPPZynG2UZlCfztWyFW273DV4l
6SdT2f1spVt2VaFj5S+Wty4UKdJvnztbe6+JYhJ939tLCW3I9rRGshH382u7qm+3k1fZC+9z3N5m
M4qBHucvhWYD6Tb2rVYX0zUgHbthtz02ku7cbNkj+KFPtCu1vsXGM35Xk5/tiMZJiAtVIYIhJY1C
XEArfgn2PusdzuLcs8KtnNMy7kIFqwHl3/fvHFVhTP0+Dznu24LbwVipDylLdALcuvm2iL6p7xT5
UbG6kOmZ+XCTf2d4gpHg1mL/0cJI1ZSvJSdU+Yl3otQiJFRC352PKaXPSgZyjvzkRYRtNb4gre24
UaSLunSw4EtluNud7ri+HST2/4zAxoXHLQxzcLRx2iSgBxK/i1qgeCCEjOnyGRmGTw+zisunXz9H
tzOstiezpopIZns2RcqmSVPlycQdp7AteEpGSIuQ7xDsczLXJpSTNTb/dsh9LzB1K92xLILE+3jz
7PR6ll+D+yK8ARC4xCoDzCA942KmvnqMFzIpl1k04PibyeIxnvq+wDICraoJZlANBPqapzLB6C0v
tMGep3tQHPNrqienbcgrrU0Gsd6ME79dNWiXDQg4pu0z0LFZveAr+c/bivjR4xhdKzzniePGKnzu
AM3Jf9/lo+ppHcDvNExRbg8x5gPU1zdejf3HlJRjQcUeON3CGAgowGPk1Q8OVpKTfIK9aaE7JBeL
1APy5SEnpSdf4XaZqaoyU45zAbCm+D7JRMKhrm1h0b6kwFyS7+TnAX7PpsOmbt2MCGrsvnHtjQe5
RA8HhFfeFWvYQKxL79txU1fL00VYGFgET/tPClCg+WrX1A6ra7r3uq/A/cYXO225QwSF3d+DLyrq
yOPpEIYtkfjye8sh5ODRXGWeBRJVYb795u1nLMnGGJa+QKHLCSwsasmNkEOz275/Y2aZ2nMoJ3NT
07z19c3kzwkWpQsSRWBMUGtJj1HimzVy9g80RuzzH4iFsxSq9BYfh3RX9+Zy47F+6bnIK35GQLpq
2/vKELeR9wYjamNRjLWlEscYX49MT1ItTever6Q904jwEJ3zwcnzwkj04FvMBqI1qHRky/v9J6mx
BlXcaQcGkqUa3r2EblITvp6ZePvv+m0f5gWPYoKSeRyHAiZZ3jevn8+S0cykEyPf+ImKOeLDiu02
n0kT6JpY9vEv8h1R1po+dzijMeGci/pGvQ4r9BbHe/jMYbQrUNYv2dou0rwfkXwnWRhGo3zzKsa0
eFPxN5damN8Ub/iBXjrjR5iSeT4TwxiCo6ufxV9pLyQjtSQA/jkBS4BJi2FWTU1u+ym6NKKszAUd
vAAjXr3bt0ME9rad4E04Cf1OLe3arSmNzYQV+GLzYhsYexW6fM5U0Huc1Z8mG1CTrpVgW50pjj1+
QDQl73dBSXO8y3zzd2gBNdQWLgByUBYtPameSRYcdBD83EtqfJxWKZ+xBk3pbq2IyfPvSkX3xE2n
VpnYTWwLbDqvxN92mBhJm7zTadhXHO6jXhcVKa6WGNgNRPycoa8YVVXL8BfHwzFOS1sKswfxWZZG
wt6lmu7e4mBVcdkxSQGL8taND/mNIbjuZJTjafoskoYi/DO65ZdGRhnoc76oKgstxVRaWclH/7dT
Nfn3hik4YZtaM1GRt4Z4wAS2vbXjoQ8ZuggAvYViT9IYrJTk/ZlehnmTMVoNxSNgdZh27NauIhL0
FdZ4TkNWJ5r8AhItR7J2RIImlTgYmuiVjLQ1hmcdpPSKJUP8dvKd8Bac1+4BL2LXkpNKqgZ6YwCm
Gnrbs6elDB5gcTZuCteb+DqFKs5Qcy8bF3o1jbuNuk6heYGT05l2LQcvTvH4+2oiQ80CTTc3Z1YX
CnfbmJb6yRqrT8G7r9jUyzWUv36v2ofWL17ZKqMck35zYZpuXx1nVSOd11/eyLdlNKGyz+Lp9cwj
oSlSc1sdCs6bL3RjPYJws9DaDaOswYiCdodMluTNpoZqIXKOrU8OB3lwBOuyr6vAsa/fL97C6tUB
X9uvF63wHY3OBAY/mQjSIDHwzloQaYLhSV9/vp0Z35SkhgzyCxjbFlet2jY0EZE2c11EJZMxbF9L
DVKHceJmVebKgmxP9WledGpXmRP5f+huAZpilUcVaJUVAd43knr6ZrKFGm2FrE4Ip7sgtFd9eTVI
V4vlzbMWzktMsRuUfhT4qYjKJMsXNNDFvprlsGZCMOOzFjYZkV76m4xOxehVfcZDJNoRlQSt3U6n
XHcatCTrWGjP1W1Lc7wmHmS/Q8hFzJIL64peF2pA1JXBGa2cc6trAhvUcl8yQuxO13Bld00vSxoc
F2bWHhWNrfnJ1Io7TTgiQU2O87cKeDBoWrX++upYTc/2EHqA4mZG8ZHiy2OwkfgqDgtUhgYy1RE3
LWqXDF/6coV9BhnPwRYqO5GXomW08PjgpR+hyFOKC7GEXT7i+Ylyfb9lWI5IgyFBgK8fSo41P2II
5dZoxkUS/0rnUwtj8Ur8+VUzWYi2kj5QiaKNQ/coIK8Vex8zYT/sCr1j3OF0aGo0IVmvsBRv1tZ5
9NQ/NKgPvT6iYXFbgTJul+B4dtg7hofGlUPIDSI9+9i21NNKmoMVHmPWrAtjwvrv3BN54Snm6/Ng
IAyCDcGvQXVReDk1nVHkC4807lJDyoxfOwr73++Rij/Ds0UtBeFCnl5/Qc0OlVzYr2v40WZBuHxF
PCHi5i5YGI66qdXf1WSXKP4vdL52l+L1jjULqfgOWJ6l+vgyBFx5e7Li0d9U6D79ERIrzRjWWQ60
LaPe1h7Y/avYOpe+37T9qFZFG5rNAToWacVVXF1Klyyrxt0h7pEgZDvcFyfwq4c6ZB4h1AsuoyJb
hTKsQ52JSeOjNGIZWYym5EYDLEe2856HJ/dfTMS93IK1fcJnZOVGdsR8D7ny4lkK06PlrjhU/dSt
du5OcM4Y2h2LM2WRxrr35L2HLBw6QVaFJgZv6uPOEJlE9kXGifEvJjoJKy4mJprkH5dC5pHGdw41
CNnjvGS4rs1Wg3Ylg1Pq9IrYW+ox5MG7R/g/o6ILN49JDCXvCx40k7bApNR3HBpV4vbuuLU20SOO
SXPPeHmhZ4W4HPkUtGaI1HsTKADbjJ8j5vW37BIihJCzGd/Z6S2Z61tvpxxiQmG76RllrdXLetO4
rjft9mHQMU9f7nRvJr/JQQ65+G099uOoES7wAGNXZD13dPtWqAXFYUU7munusdkcgoK2SOFnwCCe
WbHul+6Xt9H03cZ6/Yltpj04J/0nBvo0GEGI1+jBGjFoPT/sXJvEQFuuonLJ+6De4qnG3HAgboc2
5iiIruLLIPHzC67hIWRWuZA5BPimisZ3QRQYQJXxv5jcFH4/dfWKSXwbXFvmd/QKroCXT8yhkQrK
FiMLzp929GRWJmDVwqe0r9xFHR7cgTe/kLErDB78f5U+JmONVriCjGdbwhcU+aoYOr+ddPhohUKG
7b60/aLbCMe1z3MEztHMgtlW3kpPpF3YyNGEiAaPhmVSjFGSFIyUh4FQx6/8ttJEN8Xi2gWcyNGl
P7IAQrgNJnKRBrqZYGVRVuaya9hKdxs2dCrKk29CO/3F5YL8y9A53or2g0o2JTa4gch3k/M0LUoG
4pdiIj2767EGPqeIeAIsEFj8xsGmGjdfdIfJ4MQHLDpFSJ5dQAaOgunmjuKb0l8gCxUTXaBu2EEu
9BCvecYWFm3c95jBldPKWctQT2y9TqMg2xY2ZSyX6jlhwbMcD4poA/kPGPZULTmkZZzsAdhmBZdV
piuQ3M2NsIIoT52uFdJ5H8H7v5aC+WLqJmSnH1iY9dhH1p+XuxeV9oI8ahXJmz8tRffQ7Zw6cK45
FZ0tsRDlk0msE19N0O2aOV3E1Tx68APJcbeMet0udrxI5pRohjStcOh4hHgir+20fu8MTtEu5Wat
lrQztPwpWau1ovxStRG9hbaKbtr015JJynLew6PfQ0eWg15J4jeB5M2TBvTew1vsmcFCcMatU4p1
W0QqQzWS/IYEdfAyTf8Y68biKACtJK2nzDyVMyOvCLy8d4+VAJQih9OD0F/vBGLVZNw5V061oI/e
MyRWx7ad04Bs80NjuwF68INDhXx6WT0aRYm28agjWfAssnjbRnCNYTfGKF6tWs/mFdxa/j4w0QU0
RMNl1QfWWGCTQWtw6wsD4BEmAIFwKUvz5q9i/VrnIvUz+X3llrE2FYDkabrnD+xkNH8l+YANEdbq
ZAj5uRUAt4D3YFqcbtPZgH8mF85VRbvTnb0Vhedwgb2QwC1lRSzLRa4gkSywUY29iPcRLpq38cV8
eLKOLLoG6rw6CDOiysgjz8XsdRZr2U/+E4bBSifDHYWvol87TQxQQkrHOgM4wpz9939E1cXSDOXe
kJq+Caey7PbreSjyBfJmJfvjA1pYx9Mwf/kV6pEFiC4jNF0auWyqtkfQE3IEpOix+LXmXYQeSsy3
6cBMHDcGbUi7MFlXxLx0rGqqPPRkll1fgyr7gUDzy6Lzdx8Aw7J2FtkvLBKyc8JWFrh8nxl6/3i7
qXDSK9FU88wDCodB0mNof+4he91TGdtxzuiC1cz4wNUj3yWyRVxv2O7zNg8gYaGykHtLfdsFV4w5
elSfTi1yAbG3BJ/L9F7hfZn5jzusJ0ECopgkop/LdUs9IbnmNVXK77Ez7TpIYhTZUpmTSftzuvyP
FoIDcN4lsB3LtfIomLBwCm29gIt+6g29iIpzkCiXuWEMioNELHqTDYgruxkedU1p0R8uYYZfcHzS
ADTvmQtKU44adpbEJgqskoCNX7asiowqHSv1xoyVRPG5Uc/K0qllMMoFeSDpwltU41L2sT0Mr9Yd
qFnqDpGObDGZZXYlK2mXZot5Tc+XKn/9w9AllDDw3jppSWlvZKtRsmlX1HTT13YgjQpLfcm/UKIi
q8HxBeyUihwHjtxSkHwbmRSTOlgPKY4zu7nxdnTbQVBI4lIDeDlBe5qHTbr0MMLt7f7DDiMolZ3f
JR3CiUqhs4AJLxRVEPd7on2MAP7GEEH8bDRZ0HnSCA/9ZN1B61o07+MiMBZboRd2SoO2JRY5OPTH
hejGA0cIwgPT2Ae7mDS6uL2vMNrwH23SaLSauzCWP6G+Yd7Dur4mdicDedOzkfj72bolv+xs7kIM
UVtHEvCwLo7yoA+G30VaCvg4sXBRzHBpCbsFlTxwKIS5ORpU4/2wHAYIZO6A1TQhiH9OombhAIne
nBgCCEzNe5DlNnERPBGdkMhIgl+ujGsnDKDeYzhQ2XYlrxT8yk4r64QSdLJh3gtf1gw43Ki/dcEI
278oM42fReEGojX7cedkCpKzEMAgXIyQbgjgiIIvMtmlvLHaq235T9Sqn/4Yw+CkC6bND1Orw+Di
tJl0FOS2jj4Lll/IQAAK+7UQnK6nqAtzDBnDtTBeOCJ8csBOK9fJmkZexcyr1EbaW+6DCdZ84M6J
Q0HijQxfQ+3xbvJz+ICoqxrAbktv2HZx3Wd1pt+ktXkjF4qjc8INLwis4MO9ZvEFDbe8Xf4w/Msn
7utqlAnuqYSRolSSQE79BbF9RLCN5yl7L+fN6itUuMnDdRm9Nam2+do1ygJKjG70vNWkATDHYM4e
4NRiRCAEJFiZmZSXsSZFCL3/Aw32Uj9UpHtxSVrKNEm3KxgiafPZ5n/Xl3UDQcPDvOfrvuKQnkYy
2c+aRJwuHC6hbgygnLnP24qydC3jV4f7Orzkyj/N6uh6Qj1m3YFZxg9W/ajWBoSuqNXuRE/jHWuc
cR6OI5blnjFQZliQ+sFyZP2B6LKNcnENNYxKfrefFwStOVZsN/Smya/vEJaxDxm0/gbhEof0vTXh
Fp+MhnxjqaaSLSG9dLTUjBxUP68zIerkMf1R++/chrdW9AYfYvo/NdDp2c/+nG4FcJWQDjrIsUNT
nh/rjPniCj/dEUGCei7vjDeu5BM5BYOd9vx5jzQLheMhd9QqrAI6Lpk0KQ1DIRDmMTNB+qzcbEHl
BkVefyXWIW4POWQeJ7n+FgfBQY7akyIv6vqtVha+xpxoT2o57C67DN+rcuOPYVhriJmAhfPU+S+i
GTFBdty0zZ/O2You1YDinUMqUgzNXq51EbbJZbAXtzPyDVM7LXQ5AOeVnPWUWUu8ujoXRuMGYBec
q8/+zEtcFoZHMW+XhpHyXVYOANPqQGITu/pFv66i5QlRqJZD3SH9z4TjQeG3g68xR5ZOzYym0g5s
2mSfe3S3yznhmiZ+OeDPMyqwCdDtWCdbnfNjRXt8KVkIVhoMPQ2NM636HYUBKmKwVeH0uWyzIsXz
gcZtWuKRMWwUCRaSF2CK67+cOrLjcM/3zUJky5ePecTQke3aEd3032IpULRaKxL7vw7hmy1GTnoK
hDG4P0Jk6SsCGJnmN6t6OroQ2pUKGWGAvggqu25He/+CT59QjboF4SmYjF0k5STi6PoDZlEMc+pN
bJ1t0RccVLl8F6FRAkD6U2kzSAWZiamgGSQnhRijxManxQxivw7BqJFgOGSw2uX3E+9cjxNsdF8o
ws8wEm3tWEWaPkVyQpjz8jyXHKnaB5FMusDveqeOaozSNLisg+j30qRixBZ3YHy5PyS6vj3beV0i
bE18FyEqfxsa9sEG8PsiJrtekl1LL3OAeGvcHcyomK392T8J7IduNsj1tegahTqtB4Vgq4gFlhNv
XYmKb5M/ZeCLODhnCAW8tDFXAP+hlRPk7HGH8+E6OSoxIMM6OcUM1MfNugNifLDz9ot2vix0G2HF
OVpwqIn0+n3EMWYTVB0S5WC8kP8zToPpcpz5ulCAHD5pnBVCHJXPbf6YhMb5u5AS2YKbEQlskhQo
kB9MU9R/pKb5KP2CSuk30AhZg2hm9bx1UMputIUmhHun5X3pFE+l4H1xAQ+/58buFTi/O/LjETfY
DWPC6PlsMMjAkQt7PXURctGjmzNwffQn2xwo57+FoH4WLDaA5VFD7SKtu2f9vwywzqpO8jvrLnE7
13fjsjqWMsePPnruIJJd4zA3sX1EKguomK3oAQ6Ipj0Ru1cALAKQ5KaIqE967K6mzgbJ3WcX9fo7
zbMXH/EdD6JDCtK+ccSJd5w2Vmq6806YtAZ5nmVyRIoOzqAHJqW0cXEp4hivgmE58qjhtG4wIJq6
HKFmiEuIkvT984Q9hdZ+DGkVGZ4QSHy08kQNZQRQt2oZp6dQXDhNpEszakpv/vScIzw6r8/dL8e3
R5k2ChlTOLWrTle4qtfB2sNRnhl3S3m3beQxeF3jY1LBMN1fxvXZ9sX+L/7RxdkainI9BuRLqkk1
EusYvUKcFLSlL4moHaEHU6m4pciQ3Iohc3FAL9TS/YC+nugaFNGunT/oBfAN5CiUaK6m7q28NekI
DAFD3OSRDock22ng8ZZo8o3IIrt5rim8/mZJovCTKWyyxlb8/soUwXoAALzszH6ft96Clq34nzlW
CDoDim0fXKJOUp78seLbNg/su0MEZkHp6g+t/vbG+UwWDtiGDSnGL3JCJuoU1NE41tu+uI39rJh6
Xkg07PbHPgxtusuRVNIvlk/U+dZa4LmGbB/Jxa3bJhVZmYNw2cVbrA9QsVXH6gnV5aBBLoXblNeK
tTM70y2C9jj4746puarJNhQA1Jas/6d8+D/EDzYMI7mNYlsb1iNzd2zOwD0w/YAGZxLjVp9oqe+x
i4RhpaxaBJ9SFx/gKH1g8ouKu7koe2DajHUqT5LSYkzRNX4Wf12RHePbZdcQjeFpBotyMr7CUnW9
26QwLAf3gvhCd9xHj86zrE/CZEW+1rlejlF2Bs9aDNd1RZQa0FH50hrLgIA9R12JBIEJgHkL+vb4
nmYWiIhKoEJ5dbKfXnZi4Sk0+4rkyaI1aoT3T8yMDM8hS9SuEeGwyzz6z1+bP0eGYdZOK774irZS
YMNTq5JusZ3rtEjYkW5qxNHmvWj4AteNwi3xfGqpjSdlqwWaai4CEZkZ3XpZ/SxhlxbTI6Fi9FTU
ggFM7RTgdgAz/abliWMVeIRLii10EnN5JBahAw7Vi82B5PrbOKOjZx2G4G7YjWHEGomjw5tfG15j
i+ANviiFMkCn9kR7eTo9+NwIRiUwby4zr7bpqlb2xvQUgF6Fqx2yit/AlSV+aUkTeYklRIAUMYq2
p451JE6HQX0NUkcE5a1H6GPZY/HeIbaF4d4vVy0WmqlP7cBIs+Y8KCTp+R3Hxoe/qsHGj1TUd5tA
B4yv5xh4Bhuh0V1z4jwf8e4nOAAUTW4ZfIl0wVY4v6mJajOIA1bwmzJZUCM2TjyB41FMQ/6/LiMk
Ul5fXQ2yFJckAnuQi5mQdJKZn6t4OcIc8ZiZ9WTi+7tpAY/B9d2Jt+ZF5VE7SU20uEQEpJ9RfC2Z
SIE+ydg4/+JOp8U6ifMYt1DD8a78lpC49MKfhArxt+fAd2N5xAQGnYz07v9ipdABN93xShZxOzMS
KkktTnq9oGEZ81suHEqYIkGx9q6Uamst/+xC2G28EutbwnC9/l4SVwcR+RlfxYA3TYXeRdrAkwSi
q4LK7/T7emNQch3kHrnRn2W8As2bk+oLdFyN7UGqQu5p+Qe2gESyVbiEqDM35wMZZqxLkMv0Qwj9
Q1VaZD3UkfV3d52pxESlFfI66vwKtzH9qjfPao6SS5WCfPIPXWbVxxmnzmJBl+IvZW/bWyNLxLhe
Yt0KADPbafZiy3aB48PQipp8z4V06qRs8UFFknW3UyPSmNGKYgG0oIXB8Io31xgt6ByJ3IRUnu41
Dwzy8qHZCNC2d++kI2r4d+pV+XhpDRVoESIiP+pJ8ejzlDdq7od2p5ZD8FAp9vrsaIYasOEngUMF
HBz3dd1BXKHYvnfF7cmlisuHGgtyJWMB8N9vB71YIR04Xi+0SSfB5bflbQJS62kikz6o4Yt/HE1R
rgtdOaBK0Dn07avigGqHLG9v3CbneibcQ5Fg3QYBpxmpB/m5LimTinnKxNbWpTIaD6Mqt1RKj5QG
HIuD4yHPCsfMZkXZc2+lFRDGx7lCrS5DEVmrmqwO+6VHNXsbUDaSLD5PBX77ONh3kVGD7l5+jMLv
c6KTcdMhQE/vDnbCay9wXujXfe7dURtm9d62Ds6IjaOBlagtvcNn0LrVlLRoN4xvIGhQK6qFVNoq
Ni6vj9XcCW7faNEdLsntsVC0rD/+VrgvLxLtg/io1hcpnn81lKkC2Hi8LbBg0VSyMcvMX6b+7lPT
lcQ3IxLdFaEyFCgzANd6+unMKlm4YVtRt3ukV2JHTsHJHEnMEs5f7O9TU3FoTxVwLjfs1r/3rIZP
3jlzxUJGxPL5lmtoDC2UpD/8bn4LSuJfB0/QHb3jzS9DSci4cNePVIDW+BkVcAB7duwSOEUj16Vn
gvjcVaju+sAfDCsHt72TijdDJHxVfjrrAykGJrBRnrJ/RFKyj8fWRN1QILNI7KvY+yZUyHB5nnXV
qflK7MI9aDr40SHCUnLxzRgs3xQAfPH6Ao0FyyHUola6615RzySAXFmUl+PXKWxttgF20CxwMFIe
ud0D30KZc88olI81ywXG2AcViLj4wZ7eB/7J+JslIMMp1tS3IEeH4xUQqF2EmbUmys0Rpi1bYH7/
UJau5Pt6orXu1TeOMC2CMQIxIAJv9rOgnm3iwCj5jDCw5Oew87NHLVqKE5GwrvcvVaKviySnOTSZ
TDVcIwsutuKwQQ9FAVs8s8wcMKjtp9n84bJU/2VvQgeeHEeeD5bxe/wy2dsFFAS0z5HJT/3/tkpS
BI0VFyKwifpYj5V+OavUeT2LEVbagKzco2Tj/iVT3tO1//2kGa5fdw31Sa03oao6GD19S1NyYA4c
JHlC13O7/fMgEDTQwZPfrCy5Wk5krCH5nFIm38ZEhRl9cidn42QALciQGYUjfsDQMdMGvVF9/vH5
Obgu8xkew5ZBA/St+sZ+G4fOjdBCsl86jml2V936zzsq7BmlI4cHTTTtfz978WIgbWX0y3UHSHWp
wDW0OXz1PMDYeO/w30ma70Xc/KWQzaLzgs0/djECitkO/xXX7PKUUgfW2keCJ8slhM77YlOw0J1a
kZPc8+EHambuJVlO0awUT46top5Ds2At9F3tFkDve6r9c5Gwa0diO8xZXDLRnzSKhVon+elPQa1a
UDDCpyMPK73VkkVDFxVVxq4RDu7cIXQI4sjoBkDn61Sj8lh5w8clIECxW89pez6vx2dFcWjhd7ow
VdWhzWamkEDYx17vONwjgBZA5sbT+V+dxDJjPVNjjkfgnyQgLKKjLyvImg7/TvIv65JUCyrp2VEq
tR1cQ4UcrZvneZvTAdzTu/1GniJ+QKpNJ3gXlqu1T36Gq4PbtZxAgJHq0n6BpEmGePjBwUmqmQRI
4ddmdzIr8/18HphSPR5HTzGrqi0CLInOYoH+oTGHNWpIOyxAw5KhXqMYvdh5mKkVTAIvnVwREhQA
mYtYflVWFsrFVbsmR0kMJENL6XxhLLU7e8LIRd1LbVmApAy++3P60HRlzLMu/bOD0gBm3B0ACjNF
rtVbx+apGrwUFvN4AOSrCbWi/Gee25GHwWpr8YxChsVsEO2QezrPwyzdy93ZAYp+PYPmicR35vqo
i1FLAlTdalT29SRGwhOfb8zfTbMplf1VzM3evhI84PWZIL2J8HjLaJt5XwSpNL5kUclMXd3DwhU/
oYafDiHp04/66Uj4HPpahDWVSELtUI+NRE2KDsUUo+xgccPXAK2OL9CqzREcAI+GUyZ3ZOS/NMpY
dGC0BnISsSzw1QK0w4ia+OToXqhgEDMWAZIltq/ggPvoelmQXMXOq+Vt+ihJoSkSK4W+TPzCOQxK
5jQicyxWSfoEDJQl0YyXdyNX9u/qz0e3/Px7psBHkAUUupqAPqeAGX0lEKxdIGGbW+74ZO4x6rmL
g09YCfLtMcQhQKZr18Siid6Iha0st/9zIkOGvynSHnAz/X2VBfQVFVKwyqv8i1vhpu0yS+EBmltS
/kF/MD8P/unwsDzGUpmSHrzqcg1KAux/703FgYiRrLAAv+Dv9/baemg01VLWffNQCNoQt9kAQbgM
kpD8rlEzIDRB+62rOJQ+LQDOJf8JLrZ4F8OWWba+jQXNAvCaVsbq2Plyk3pLCgmZCOZedLaZg5JD
sOalc5LA4p1qFBgA/Pz6JfdLArLe729hcFClmsFTAJ3TjIdmS/dd36o1PvmqCeSazqB5qfehA8Et
SgBhE+g0dOUE6UZq4Y4yw1/3MuSGAe01WZtVbMs6QRWZH77pOHFilB65z2nQQJfFIy29YzFJhZ2l
wEHrtakRRpTWMm0hxnaa4Q8YPCZ7D1vhmL2Wi8+FiwqV5eRwuvANpnZKJgnkutV4/aRoX07QLt/3
OFtfXVlzsjlR6Iz+BMep4gVu8a2VwJvgNo0jKbB583fmyPgFlFQbXh+Tq1aKhSvbBUGb2tKqbMt3
2BGUN0lnx04ErpQqGSQMdB/CkCtW8RZZrGa+XmDuDnw8e8ZzvMTKTpWJdi5MYAX+P4s3pQyg1W1f
2CXBefGYTyt5y9ZHdWkRButygbhmb6tDyfyqgPSdzjHqFk0J2660LKX5u6gWBaNraBzAfEB3dSm3
Q9/k1Kbn2RU3Pz9PVq+CrGPeYU7TeRCgEK5FvsQmGTBCLnBxDK7MYgdKFZTkCjBf1x/YJDhJVZG9
WeF+zj/S5IWVo058imAeKZUi7HAL2GYWO3bIUlNVcB6mfI8OrOoCVKd5tUBk3X+zN5XMeGrv/naJ
MBKhH7lIH3xfjzUsYmxmttJEAjy+AHAfeYvolPiXhtpRVAMIowylMqxvXnrm9w60mbwVpWgD1Vec
3EyP3mejWIY/nUs9U3Or/M/B7IUS2nuJrA5GnqwlHejf+D9Zh7BzviPW/e4sQ4uvpnJUaj3zmuiG
5dJIYrjORnxltGJxdGJ6zwwvHRom47nkXWkoRImqDRdLQ9bMTAgygNC6l9mPSt7x5KV1YrNymrrX
mcEUWCmjiEIokQnBf7ey/Gs6lm6TFk6ts3z25/jM+TnM9G6xqjI0WeSBSw8Tiyz1D9gOaXmQsHGr
qTcjpPWjyRYT9sUXWA2/jNTIC9IeiRMmf+0zsTAZx2GUn3Yu+vsEF2bI8SD/QzDjeU1Z/6dFEf7l
kQCDrN6R/kUeF4KlO7o0gHL8zjLfxMk4JSvSVBBfT95SCkLt102vfJW2sdubBEgYyEB+Jbya41hU
cn6F+moZGI7yNuAldoH5vvhLSC7wdSMRDDSnvBYZc2OKc4gQgPXFYL7qVuLDKNR7zeof/IwApL95
yJAa+FPaEFSyxhVcXD8I84vFvQBP4jc1i+unlVMZUYUeCL6ymOxWTroO6oIud/bDWlyiZPtBMhRw
hiim7kVPWkDjP0hk9pTBPVnwR3sRQluk/kKu6qHpJPGEWH5Lox0mhYPGNOA0S224TVVVvDsFqokV
mbHb+S678bVAKgiXxmekCe7yyU+cN9vA4ut8AhIg5wdDedN/nUSwy9OQ4UktoyYlxceM6MPkrxXU
ZqPwAcBh6VDH2O2AXLiXcIwAVLXpSfApsBIEygHbCx5vJzTx7qagFyz/2XqUfQEsNvuyuwWov6b4
OS8J8ivr5vcx/gmIdNQptLSp8KXjk7jXnef+uiMiDwe040/8MnWKuMmjcqMv2Z7kwNxIA/kZCXxy
AJT91+jAEOZ8Uy8rwGRJBzGIW8CLyvZqdKZXuJkp6MULVQWWplK4aKX+7FJWUQog/1A7smKzhFY4
W20TAlZyBxn4uzcbfeNchojGYzT9j9q9YLGgZ80WPPffV2KzWQOLCAsOIvzw4bTxMRssC0n/eN/p
JeWu8/Rg4vKwVC/W9GvHeGcy2DfAZoRoQozHOEEa+NCmOs3v1rY7+52hb7TXSn7KjAth/XJbngrS
g+PKyVgj9LJ9QM0qjAXiZ30ToUeTQGQFqfeadOxaOZbqkJj4Poa0e7fGpL0roGiiGPc27Ld7Z0/W
x9JxVe1dCdmYpYaz8NMtFjQz522OegnTBYsPrJGggjvmBetuV8G79D/zrZKLO5dU5M7KalL66DMH
IyWzHcqwnvWhiNnCOplaGsxSEGGeDnRXcmWVXWoMXLgCQ0PjqG2v1zcC5TYoqk/luDSbsomLsqJh
9et6n/RrDuaVhgyKwBVm9BVICTTI4+HoaSqU/yhMsPI36i9HSkHsIRbuQCn4CHBuDDkKiqx3ilhZ
KM82wr1toOze6OFG66cmdgT335vjlkC9lDuYGCJZmgFebz4081MhqNjosG02o47RsBHmZuGIVe0R
o1Gt0gorIhxyiPpLgatj5N2FYmutmzR+5cxbEgVEfgbSqNiJAixraffKVEl/ueBlBo6tikvekEAW
E+TZhzbll4X3P/w7Pl+UVfDUt9hFEnBFNEcqWYBB84gWtRhpbrnZckqJ9x/cnFBJnOd5VeyXJvEX
XNKnZEBFGfhZKXoAe83fznXZxGaDtu5bbpYGALBxgxY41Kru66XfAfCmUhivseU4bdiPC6P3p9qb
fgNvrvEZx6dblMRgiPxq1CZlLIK1s3sjA5McC/2Ke0lteDuZxItF9wP0Q0tMQ5cgsCEpnGa5gxus
GgmE5tpY59HqRNb2CpPBa/erxFjDu92HJ1gH/sJnWuMzq2uZhSG824xD4XENi2BwzSpNnT9rIspo
M6AD+PqkzguCRVxh0WHxr4ieqg+kGyEDY9xOGmy8Ol6bIMRRRNRj9bw+SLvoQeu58Y+bR153bXYi
VBzJd9xKXn67sLrZmdjpa4fiL8dMB08jOWWfWNAfrl09VvAaRELKsV9X8pE1TeROs8X9+haUkKnt
eQaLIkVGiVr7AKMXjM2mCBKCKV+Yo22DQIySUGSEH2wxokw63pWK71MgTkA3NDmUUbbj7UazgsO9
I2gi49rdetrLCXRSPUYRUOvDna9nS2ScWWLT+xj3zt7dfX4LWrtW1rSvqMzEH0cHTENPYZ05UkcI
FKeE1YRQfEMGlcbycqRS4+83IKHe6yn3a8qR3fxMbnIkCCLr62THF/A8mzDCSH6uq5TWijM4kVM4
YvARAFWfJ9AWxPb8leM5JZKf8c645iQyuAd4FW0HQPAMxy6c7uZBtNHTu+mHEpy+Hd8MB+2ugfXF
U43yuKzZ4dfU01zl6LNEvabBm9GbfQ8tBpXkgN6s9yGcfju03cPlr+B6sDyHcZfpHchlK/7xRnXD
UXu6DQKRuEYQr69FKIVY13i5/IOFJG0SEU6Twp9ZdMrjL9gUKSC05yTJnfkADwMg3PSMjLndIm/O
6iiKOjRCJgN+yseIEe+WhWwWaDC3hL8W38YmQFGFj1thWOujnHF8Y8DAWlAHRqdcrB3PfonpzMf1
uOWpADVrv/NqRsU+N9/BySU8oED5DwFMQXujo8NbJA7ZEyd1iyCx2a8GvwtIafW0rjqVk5O0JjO6
pde1vblCVe44rngTBdgLkEmL5Dt7pDA7NC6Ps07BZ6TPSOqdRn3WX65IbqMyhKjKaKONQVtqCC0V
tzK7F06BdQHZfJ8DN5i45JhMUmfSS5Lj6gcpjRDxEwCfMF8OYRuOrtc2jEzpOHK8BFB+HEFujyb+
rBTZPo08dmyXL/EH8qKVxTO/VVIlrp4aUTP48kpHXfEDDF+lNL18uAUxLFRdG/yEeCmrQRF6DC8P
FbPhLzGiHVChnw3sPCfX6MEoZhLZk2SgyMr6GL2tMFo7/qYNvENqvSnmHoKl62mugLQ6BKJx7j/w
hUXSt1uPVwgmhTv6nEV3RUK1nO/9t5Z9w0qBQ49vlhV2UKTJ4Yel8c9okN/UjvnmPDrInvUFIVH/
lqqSRQ8SXsGaj4kh+djfZoApRMizMHJCBNH73rntghgqRHaY+nDoH9K52zjnkowTFnIM8odnMmOo
0WDDhR9oxMvMb/y+0HGd9Au6rxlKfAXR+Zpr4ruz3ZzPfLlONPWrtOYyrmG/wPiV++CJds337plt
16sG6H0Y6nANzwJyBcaOXx2J8sdti53qDkaVeyXmV9hJ3MqjhLG7upUf/b4djKxVTRITp3HIELab
eM8gxOqS/y1OMh/MbrLJ4y+PynvcYUDlODYalyq1n0iBCEiIiHQhjMKaU2Q7/np35mCN+TOVMz7d
yuWu11MTOuWyrfctWGCgHI2yU9K1nmmkLKrzjdttra1ynLWQXZov2oP//VZBGDma92hZT2B4U6ox
ITMGlZ9jc2qD+q1QTlmSWN21isM9nWDGz6TIuPlNRbXWR//2aWYMOLPozjLWSsmrb93OwC1qVGCQ
iR4KlAGmTsEsblU3tcp+4/LZ0JZMaCXfqa0QMRFOInxuU0qqCix/N4sQFjRIJkTn5f5raa7B/d6O
zPqdt6iboRTnckzmToEjNqU8qb8Bc6V89JdgzAllbW+3fjOuY1RZM+IzmQnFxfpbYBrYAOFdQcTw
3ozTs8oZ8YcJI/jIJt7Z6eGjHI6W11wos/tx8dbKt7wFWaD05Zl1SPcw3zaJ+zT+6eOd1f+kWoST
kJUjUUs7ytjSPSfy0W05S2DCfgpZZQCHx6eRFnvbTSKDlIXblDLr5TK8myRPUVUXgZKiUXrPMA/o
yY485vQDctQd61hhC0JjrhMf/cetzwkCAM71FM2Wu/6UGginFgdOjpkm/XXSN/RaxXDwjoFlxX7v
co11mXrY1vacPBlzqT9kXXGJLvrRgnVZDTj2slWCpnO3Fd8tVYa8DwLfbPjn14P4D463KP/2evb/
LPKLRB0jC5FXdivtkiuYE0OGEjSt8oftD5xkXW7cCDaEP4B7PtuGh1b9aORUGi7cxu6O/DzQRsh8
eAeFyTANg7/I+f3USupjXo+cjpOMk2nisR18FxU1e8i6epX/1/h7vYF79Af0NotngoI1P+5A7p4v
bEbw/3zc3HpK2pcuSkTBtcSY5+UFOFdaTqadH42ToCfi2Y/9DA/V+oLv8Lkwr7TdlUCYcRRQjEeF
S2/nEKK8mzUISRhRo7wbKlSJInw9lFtNV1DkQf3+kyH2f49RCuQoXgkxxfyiy12sxZqFy25bZh7Y
S++gaBFlgsFo4MYgRUtHS0xKO4rfML3HcFjPRbJbqjUyFptR6DL6bK75lg8AU1SGVAviuDyuZ5LR
r/N1eSt30dNqjNub9Wx+7qTKL04Z3EhxWpK+mKH9xA6Q7XwVp++hdBz/1SnyKex5NfSC+jYZSmmA
veQfYzKxNHR2nifGzbDlqlsc8tS+Iqm0dimPenoMHdaWE8T+cp+G78xZUYcQjQwrRbzI6cGUXr5Q
LcjuxMz2PaUzScKyLGdcGN6EDAREb42VI7kMaJ40Vvh+DIbSduXqVk2//ub5U6PVZ4vDktCqx0TH
l3qUxpKDr70oiRIMlYYPe7AK1AE/IT2oEeH9Qt50yVRoAWs9CPhIyf78/k93n63FNg00d6h4cctf
Ekk+zuSLt8eGWjiC2BziPc7jWUAFSH0IRD6ma8DK0R+sfOT/71Xao+KEx5l9NvOYKUmIX/CHF4Ps
/EDt4tof3Txe01nz6YykfR94JH7SHAb9D6EOIv8B62gFv6olVP312ZOvaA9eNJKpdDUGwtpj8Krb
IZ1dIjlBuQ7gBWlr0KpwSmVfvMzzfHq4MQviMZVxh3xd13qmt6nH0Kp4pnsEwwZ7JjfAw+lLyciQ
5NMnwVgA3D0wdo7YZeZlb2Ny577lhZINGHp75huGVrhCzwmmcIdnpsaQ/SKPFsnfCYHaMG53rgu4
WloQV+tc1RVa5fTLtKBASHoViL+U6Fizn/QsvArU9VhG0BZoDDpN9vWcVoXliUMC8FcGoky0a0GK
rAOEEWmLgXjDPx+axR+pldT6eeCR0lHV8sawBQEpqyOLviE620fnIKC9D+rGpGHmFELaePzbHORo
ZweQ7l3aZeGYpbHnGTsI7KPAha6s3epb4bFbCF2jPrlumPwzk1LPBm/FxuZJAyNkMMS7jK45V8pu
OuJ6wDeOjjfCiZ6hggHO8UpNb8v1auBE4Vu/4OF8/QR+SJqS2gEEy1J/37qsYVcWsrLo685alpMg
iQGJzAKy3S8NA1zSSwZK/gnqjX9Ae1GXBV0fAA1a8VEs76MBpqGBcnzVvcvNRSMkKkMHPTQLW+A0
Xrlk3XfeES6ZrHNJCdnz2QtdrVBRpzzeYM/JEGKEqSk0bGPJFkafVcOxp3gwHI02v+d5lwU+w+nr
PxKyPbn6FjLlH0bRuViQVJcVsb1n+zeTySJPFCbIIKKi278ABovVew14dY5Oi9YxpuhItiV3PG5C
2ji/NeVWUCLBhWXjBfpYk3MEuypPc9Hzx+Ub5x+hWo3ECxeyf5DY1VcNF+2dKtK649+JNT+VVYMm
Ah591lNPHB1oNEpb3wps5dJYeFrT0OpNsMA21biN+HwwPrU/tRCqgesOZ6NpIcS5nUu9VSLQ/HTy
h5jZe+6DXp0wCTFgXIdChyNOMC0v2cUgSDfmomyD6ekLa239UeP0tw3x4dTBG/xq1hNaT4h8dVid
rhW2duimuBBiWWvnLbq9NtimDwRApLUZ2RXnzm1UAJsJkVBiSZAljRMNbCTKQ9y5vvVf2t1l7Xm0
WyoEkvC9BRtrGVMX+zVtxSTYJKYD7tA0i1ONZfFJPvL0krQZR1+WMDJhBWVc/86Jna2qnyb8dhEK
jVyKIOzFvklOsx4F+SXKJ9TTlbMF5PpJ5IikZsVBn1d9KliRqI+ih3eXt2x/clBVXlmHv64M2ABv
NKJPjokvmVUEGnldvzhaDa1uVnhFL3KhUHkR/MZrTFKg5z3iBhO/Gdqsrg7uELWEN1IENJqEgSFp
qAuWm60/sZ2lbIDQ85aKBuwyPAz1EdUIOacSQCBgn4w7LYRVqR2gd7R/xh7UuhWyCEP6Q5/xSYL/
wnL08oGIPCSmkADVkcP/wn1s+C78gRKGJW7L0tfqySfNKSwvtLD+PzjCygEX2LLxl1ojlgAH0rKV
6QBl4c0y+ATvm2mjoDhOlGfFdQjkps1U5Sxo6FKL2pYdTL9rnWvKfyelhSTlVsOIENx1z/6z/iIn
pU+z1DiQ8DJmQVQoIDV4t+yXPTNRDydIt4SCPhnEIPEXFalV+r0jUyNHVEedmC9xlWMppFpJn93t
Qf89NHVS7tXealiQuqWRasLmJz7Rpf6qBhMDW7HGuEZ/3QCfHwMF3pQ37mzi6X6UxdfmaYljqAX7
caJcPVX+iRhWnfucPu20ipcXO+Aewi3fmMWeuu8FtIepmsPneGhYJFkGaNng5k0T3rg/StrJGRx5
iuElK6Ge4hUaRA/TeO8MOV3ESqMgRPcxCHT4L3FgJ1QOwnEAnfcHESYoE+JzMxAgsCVoPqfhOKzy
jEY8D70A55R41d+TjrhAt1K+C6Tfo9osoTMvTtUxEO6nMSwFx8lLOkScIh+TDl4hdwsrFueRTLXi
AMgcM6afloxwMkbFOCqcCrd2PUVeRPDznSHXYghF4vFS8555oOIHM9TPHi198iLQiFCoGYKHTVy5
I6L8cv9zJNXJj0atiP6idaN9cZVVwIJZVuB7tJVCSsZXWtgkb7/yxqfhNvYUtZkiXHN2QmDkTvFJ
1bcQffDf5aIl/XlmOCNyisdCLkDT4a+4tmY09DZlxJtBJFSsHh0ix2bdLNMi0bh3EvTfXFh/t0SK
QTjjGS+DCPAnuTi6H/B+lv0i61ZYoplN3XRO9vXzqqAplFCAGcagDOZfMDR6+QvlBnTglYjdjLkJ
Cnx47sSTdR9v9Hija7OYY32mlr7E7Gkop1Kp41oHeuhaxZTq50OTGPkGM0OjcZedZ9KMuI2ON3pL
dcLkK49IL1ncIAhSne9U2dxa4Y5a625+UQstqkl4IKRZt9i+meVzekwIcYernVhME6egMfkKxDhE
1D3HLBCNPjKc8oOEJHmthYzh9WlMUGKzYphjRy/b+kOzExdDRdWIWZoYSsnM7RA120I86jtEowH9
8+0JS7qLKO1lHKtydAUlVexO/SrPilxTS3g6KvXbQORKs+V1Sd96i6wjCGLHm1k/khnt1LKpqr3k
O73mvxsboPzqlB0yBr3rcNXFQ9k/9vC4pwSdssAJB0FVKDzvkUvRvNojCGeMIFhsQjtE2qniElKl
PGFVEvwZDuwENhpB7NsLJFsgC713mAo2wGyO7VFT6/In2ytqHUzJkfsaz/hUvN30uuKkQ/MGlpE3
zSnkdqZ899PBV/ssCNh9DGf55QY8GUiE5IsA8WLwd+NbWQKFH9qRLh5ZvrXU6c8mVPZ6yPknPIxw
OAqFKQgn8tjgjQY8XGvi1eFjVKg23y633PrnCVAew/cPBJ8WAHijUULNrALu39ykTS8vpIDEtT2e
V9WfkfF62rZEGz8HiVlHeysuQLHAPh0kOtQ95XBk98vuNxjH0ut8EdZLd849R2qqrGBi0Sl7RYtn
R3hwo+yTwl1vu7chP72ODZ78XJdyZc0H5rEuiFHqMs8wxTSI7gfCTLglDEa4qLipmb6fwG9c5Cvf
bvcu2v0LcIK24PdmcMPeEJQuPx0WplYwStmyFb63VBcdrX0nfJY+cKxSAIQzg08oXqerly7H9HMH
SiLRiOe7vOwA8cJBIDY/cgt2O/tlOizHtd5ETeSHOnFq2MRwcOcNtasp6NK5takLae9/WBJ7rF7O
qmG6HE28V0Ubg8Ju+gmIzBuQkK7XDysiwp7jfIHcwEz0GsAvDBEyLCtuHTnSUU1KgMQ0YKcEGThG
TRxMIBBVCk8fiscs/OkBtrmkZ/hFL913s7wEBwX5sgysxFeAt0rVOF8afDif5z2wJmErr1LCCKc6
My1kYJhN0sMoaygsjk2UKb+oXnSf57hYGN1xAqrJ75VhU5G1nsumJaa+S2SIgS4rR4xpYA6BSX40
XCWU7YR+5e9sVztrbuS4AHFLiUlq4mmorjh/GFlKOeBZ/5je3HW1W20zC9S8vL/G/OCnKmocgUPS
jdot8Dtk2mpqMXy/Lw/0XUahIl3odvMzZUZ1jxwApFFb85XSm5zKiLYm1O4bmh4K8YqX+aZcnPUG
mrPCC+Yr0C2SEuLRR9UsEhHzxOOS4F4NU8yP7mzD+uVZJR+fX6Kf5r/B6a+37Dyru5XPEC6rdxjN
3YenrLARxEsZCVdqyMOM6oOx5924RWA5g/GZ2IPEvgZ2RwxT73Xm6sJe8oWzg3C3GqwVI996Gz7I
0Ip6ViO6PKtyQvVAZ/VgMfUcrCREH9iLRICbgU9bw0hhFZBBSA4EyXVmjP6B8NpMGZWKAer9fRaP
fslbvFM4BjC0K1syErQEPanf8KWJIuDptM3NmOMs5L4pyuw8syX/mx7lVOBhVyAIB1PQJaDzAba3
Y/nMKOOWFeRic5b9QdZ72vLXr7MF7/54UP5EZstENEFvwGVJ5IVQQ+BqWRewzT1HdAlA4lQXRLu+
kXSay8zE9f6dydb8fF5BhAjI4amNyVVpIovyG8tyu32x5mZJX8mBKanCnAv7c4F+Eaja2Y5gfad+
TV5/9d6ez+1OEjnQ0CEs1sF5hJbGYCQxWBHagPZPl3Q6rZyB+TeVbUIJhM3oW99Y7/0mkn/4EsLO
61D1EbKsZDRryFArW6uY9c9Ah1xWVp4R3lNoFwEsdsz++A2f34ctDHpYe5ayBsNnXKzB3K2ze+se
Za7tJvyVdhqNZY+Tkcm6j8OAWFdM5bA+Xn+ujLCfvVgmgyI616fneOksQqdPp0igdPtPixb0KDr1
/HTKZl0VcBkseHNRYbgJmN1Mh0lhDN+07rXeVj6N+LWw4e9gVK3bVgDF/mPuggBPnP2gmB2wi8bE
dcxJRrPV7mVtMwmm219hwtF72bbiVCDOe9xguhcbkMKoW/pednZ8iLzsfJDwWtiGo9ujnTLgbNsN
Oqa2G9LO3nb/kur2sdA0fxwmOkxqy78VveMPXgmAMNRZq+zDO5kZghI5qEn7J/X7Lh4dOD9so3Rc
3R1yQTeq1nLDtyshoo0SudTmFIaENe13W+tpwnjKh5b/sGCMieh0kbe1zZO/qaJHHu4vdJ+xPb17
7aVC9Y1w86JE9/jHLiq+kMUmTw11FI09/HbYZjna7/XsUOrd8nqHNpI1+XJCa4/VCPR+AVCGc3R6
nMf8kX7ddnvQNJ+JIRT3AVDtk9fgVKKwPARMiJwOLtbFCCFvyrI1CYCw2GyZouTmkLUIeiSAlwXk
k6YiNr1cNEa9Md2FuK/7rGJS9X42mwiLmDUIGdUjNR41S5a6+GBcJiqXbOeW8pXuXoWh3+riY16Q
o+n3IoFI74JRCWdGq5RXQJsahf8jb2+1kr3ICLJ9/vHy25BCk5Hz0Jv8WvtdKlnbK2Q5+T0vE+qL
uXHUWyb2uIPElyuPOTazj7RJeCwYZUJh/JarnlP0z+J/R18XeiNrqNOeASStz4m00CoklSmfPfW0
cbwQm+R0XP9c3JZHgf1kbhXZuJfGd+9hyXqDFrr+IlXak0o/V59BK0YC+mIrRbv14tfNRyV5NNCQ
pt7uNz0xI7YquPXhtBajJiE5cI3xAoXgNOHj+q7yy7b4GaXzuF4PqpVarNirOMf1UJk0qBcL3PGj
j58ZMl91zvLMKprYHhGoQC9mgqNMeWZ3yaClwFSSNKLAeOdDeL6rOXEWrXiGPGIS6glS9xzAAnOc
jwErscsk06V4qsDIXymhf385EF8bwbdjiLUuezec/2CXH1CGf5LFX3jhrfZsNGak0VPXN9+mMC5Z
h/MAZ/trhF31bBUD/dqGHVwRc+bLk5kBawYzGkbMRaJvmGybeeEDPY2ZVmlactBrcR9wTD7+3AJ0
RKMC/1KnPO2iR80tJafndyV8fdJv5jULqpc6g4o1oNzVh770F7g5U3RCSRRjrQRHjwkjln5xL02W
LRsKiblJEzbnlwQOFdTma3+XARmyHX/umpC5E5ttcywueq353nZYVFqDh1bz4rhbRh9Y7H/MyxF2
pWxsstNe8m73F2BYBdUe8bWRmqbxbT+SO7NDMMZ+stsSZ2dApRiZO5nuLWCmWHP81Phf28GkjcSA
hSWCdO/ahIlK9juvie9F+HsPP0lzK4rp9H6OnxstAYhc8KQMD02yVVQ0BBzkhsGV9lPB9SLdpBVV
HUBr+f+jUfQOgxbd9O1xqOaTe9e9+YI9V3FSfewr07MX+TCAxx/07D/XBlXBchQQsebF6sSlZJ+2
wH8xyX4Ck4wkjuJzvilnDWHlDrVvfadPyg+36ZPm4xRWHjLQNmDySgWVs8xBphBLuk7Djs/d6dy+
hiyMkWDsEIx6779iuAlfoFbk8JUsKUFvGZKFFmHMvDn8d08V2B5P292iXYvMJ55HJtZckNfKQ2WD
EukEsUUPxiPMgVVolSUBzXjWai0kwURUA8Az6ebpz4SFkUMwwpqzdgJiuyiQsEMWuuhNI0iAuQPU
TjLJEWEB5UPvbAKDAOBx1wc0JZxwRFgSJk82r1aVoZQZ2Dv7qqmi/yOG6JCadcWUulZ3UeLYumya
+dcEr8QkJi4si1jCWQLZl8bddfx393jmqCnat6w88E7dt2e3BxwvnGzFSgetTO7KZpeHNQghhEPW
BvGv+L7jD/XNPqg64MsQNIb+98zRgkViNL9ulht52N4E3QI4ib1u8dCDCIGuTQb6Z8wUIX+Sg139
DF0KCJT1kDpJXBj0rDmM4R6mZWK6IpvTgkx93YmkZhQfhULVm89Q5ppVIIKJADIk6hntyoJXezsC
VPXmSLcjVNbN6DH84BLFmqbdIPBReLG4MvHV77RW9weUsyz9hrlZhSZT6CUiR8Zp4kIZ4nL3paAb
OV8dppKYV5qhFY2wk32gClH1kFS4CMZcWZE5a0INZfkyovZgtlt5xsxXz3OFhtWNw33U1FjNGzHA
sGVfe0Xudo2YsJOOW4QDZTzWLC2wHkMUJ6OfH9gCrSW8QxnzaVC8DukNZixgSgSJk0LMr/rdne+l
3NueZCJpVtXBzcOogjsKjSVA80sXfw6uOKjwm9zrbtA0XO6niByylNlfrN8sniwTLKu+2f3wCBW6
f32gT2dTMpw0Yzk2EGA6gQYyjzS+reh9KG9qaNmhpnDfmYJKjxoy/9StrP2nhtj9JMONf53WJOeg
uDuMIBZynnqvpn9Dhv3dqRhp6TI6x7it1TlxfTtTw18ornPE/tK3YIOfYxvln4cARhrlWmy+X5IS
2eUc3E4E3Gu+/r8cK4jFmGbcolLTl+aWqwPaP3Cc9/m3BQiLDeyXlU6+gnA3ph+Ha7F/qQBQkCUd
xYiL1E1d3qobpDlDmC2wUGm/r3vKX2Sn04r2K1LBWWN+nk1FU4KYTXta6SR8nTIUbaZKWbrBqyL2
LoLj1Ls8mOKo9MEFzA4cbtRxAYwyryFBSdqNzTbWchpSzRCXbM+MLdviilS/5HGMjM1YIUL/WBuT
vu/O+RPtrPqTfhY4D6UTmrYQFlqA6OrO6p9pQI3qpLOA0iVUn6yBN9WaViVY/l6Rs/yL3aBb5XwC
Fnp7T7zRnIxIoYgodV4bLusxLTpXIcWWYb1tV0kdJkMnXbU//yx/YtXMwp46kOGDlcuv6XEDjHSr
cQUkBV6fptP4fJ1Kf6mWYo1z7rc1i3qbdfic5JY0CircpxL83kGtuFGcI0uiVlmTUoaUwG5sgGTq
dcO3XrcuCBsk89AKX0PXodDqdoJPr6UgsJSzJ3Sf+wfPqQrTx2T8WKDVTp+i2i/Y0ueM9M4lef5l
tq5YrnN43MC/GGhLz09MMLQ3hATxLRgNQT0DdrIIUoQPWp3okmH7WD35uND8iQxupFqqOEW57Gxz
mxkyy2x+eO0J1ixM3J5BQWuC6NVLhqyNbyQ7VBYwNxfMhwZ8Iix+4rDUL98xVwgT5LKA1WErZCEN
dcce7C5BcSC1bP/GkLJiAJL0kaEQVcaxx/vBsxOnDy37GANrUbwVJ55VJDZNgRdAqL9EjXggTl4M
63s8CrBfJBvxkslq0hcl4P96bEYXiCUBpT2xEl2Q8xqDi7LknYo79Z1YVpmENyKOyMMxj6KvmaVR
kekT1kAxgpb75hR05Br6Q3nleN9qONRjNVRcX1CBECfs4Iu3NsrbajM5Xu7iWT+Mt4Yqm354W6du
q+cKF1iyq3R6iBRT3k/7KYWAyvh2hKldwPiDcQYPIdQj6mlY6P5xNrzJhCG+2rjCBAEbcZ03ILDJ
RNMhcYlB9DUxMqtB/NpmY1CBrE3kH2gTgriQo1sHEwEkNt2f/E1zOhzpAIHKBS7Xzk7aiap57fqL
qVxJx/FSOKYbM1EDkZRpT1RvMyGfAUm2uUBOacVLKQNrSze9WJRG8sGWMwU6rk6QojZmCpfAFSTC
mxmidJU9CbTo56vXPf6QKhD7njVJ4yQAylNrOTnVvmdpgpkuILp2AIPRpewJ3p2oFTNZUcOG+lwZ
hT00fr4JNQsxHiQeoNMqoUPBaFyBlHYT7awlKOYxtESW7i9QZrjQUozNSZNuGZrxyxyXOcFS0mMd
KN6hh2ces/vBkXg0GgeU3ddA+Vj2YfmpmVf80i8IrIRBTvpjsOvBQdlI/iCWlyTHmccnsja17YFe
jO0rT6Aq/JhY9fhnRHcOwGkABf4r7hDQlWhBgNs02JdmyGJ9xEQJgbI3uyrg14sDlA8L45osVuDL
4QXbZXFtzFk29jC2qGRpvVTZQicGRa6FSYs13PIRXbrsWNULUn25D8BmVxomwnEDvM0BmRuGfJEp
xJBV4Zt9OQkihlTBpLpg6e3+1yIYfX4VP6J59OF+yFZVgn08bCGytdkka+Awl2szHSvzzeEucUHm
WkZHmVhLi+OyKRfBA8CzfOcYNJCfPAN0HSiKArl1VmYON9ESOnCcSbeCccyvt+TQEx9n7ClizsPl
NBlcC9WkrEICKwN4Hqv7gPbPXDWQ6axp4K2aGoXV2alBYm2DfvJYwXLWLuJ1fLy1ERhNMOaGjMym
RCjMnd+6mEFQVgaJhL81ifyajYutHcAaAEhNtVGF8YMSYBani3+I9hqN8gnd/YM6wl931ZYsqdQd
px3D4yfNk1f55UZaD8V8x/d9xnzFXQuve2kXmQdKEWk8WJ7zp+QX3drmhqd/VPbUGg0J7F0JHrjh
F53wyIPr5I+l4brt2wRJ9JowKIa1oDzLDLolUmQx5W+/42Bmw7vaG+5D/6IGpW6v/ElEC9wGFhv9
wFQQ/yJPwbOf9lcKv+b5Mukws8sB6oZWR1qxJTyxIjq7/pGSN3Fnim2y6Lz1lXgWWwRU9zYEj9Un
/AZPnFA42Goia9wXpWFQcE6sVzucbptWFIFx0X1DhRluC5eMgmj1t+qPcQKRX844Y8PKUArDWgG/
8W+cLqub2hEn4vUTj2fGDC1BHqReaj3ChrlpdyF4W2i1aevgJCsgRyGToh0lH927dwEZdieeOa5j
7ZJCsqeid/erZLzGo/TAc2luh1+hirBb7/zVCkY2UXzfrp/1PuE+zL4ZfoojpXSAAvNTnuivgpQf
ovtxwpbPJ5Pz56Lk5eldGzoQT3zLjbVg+7cChrPAZZNMb4mPXrrIETDiGqoRPCQ8x7oOnzjPv9o2
BIW4tFwCPblaaOFX8WOuCsluBCE4whJqH2sZwX/6hKMQo0qlBPIeUfZ/clZbxJZbAla3Dh+8N0di
LCgJwRPqUnNFzY87QqvqLmjPhpbfIjpbVZwyFt1wF8iY9/YipoN0OKawNfLwIeTnaFPebdKD8JPN
rwCWPGtnf3YnS5LfSyhKgqbzi4xzM00yTfWi/k4Olj5tvWmvQFrCSVvAOsRLW1VQWYoxiId6V2Ll
e3zfuGGTJygqFTu+A78JOT3Psz3dgsX9V1eeCtNufktegWnxTyLQZH2ND+pFh0XCxkqjO7SBtJr0
BRTG7XQg+uTjP15Cp+j469+7At9M99EPC8nmDDRSDs4atfMLG6m9gtZ9KI9fT9GU/9B+QhEJtYjB
abE1g8o2ITxhsTQx4JRRkW+w8hbQh1l9Lc0zquG8k9MZxBJPxgGjsENfDMsEANiUCbAeaRIAQJec
hz0c7EkXWVeRW+3tyz2KwESPKnPY6dU2W3gyXIVi1PVrVq1XJZRwlbSeLeQFnzDosoAf6sSBnZnC
hqSLram1m441yZ+WhaamlKJQ7+jj9bvw0c8py8mAnX8wL2igOHqiH8xChsg07OCCOILflNtGczP9
AJXQb36OvtMhVePOjLRYc2k+Lx0ol+k/O30WpyzUCh0lBLMVKngrbSTN1hwG3TIVS4OW7r4tSOqC
eZLdTeEDLkdB8h8xw/s1JD6x6h8ZyrtTB5uprJVxhunG0J1fB7tbOSa1q8r6wMjl9H48QKco1C8e
usISnanwb7bHfCSPTkIDLxzSZrjUxBtgzXIPCnkvf4Z+8VvMUCFWRe/w/OY9m7app1hv7ADZyN+t
mOzAJ8SS0ubLZ3PVA/bRFeygS8n0kG6XrGifzAbQMxO4Ix7xCw8aqJdJeqDsHgiGx+Y32Hk8IFbI
iazER8Ao7mTkN8YmaAk+lUvvYfInRv2Tci1w5mRx8h1/f5XxxonIs7O7V5kZgHZkeWxyOhfaUFmv
z5TRGanyDh5TPrSUXCW/tURcfy1sDaViug1x7zoAfL00sDMq/S/qubgCQkUkeEvPO5G3/lJCtHvz
UGvoFOVLqzGQwJfc/vFEJN6thAOyoEuBhxnUcbA7oQGv3ceMMeZIz5EErR2f8jCW1H+5bsrNDbCk
8sKfKKGps3+uBm+kX639Iu1yRUtZlWz2BXnzQwCErm74xlo7q3YGDE0e3e+rsblBnArkFtLlFzHd
Fz2k8Cw/1ZIzxcYleSgvVKEWtQXWFq27eZ4GAZftCJWR1ar1wB+dd2KfqqYzfTzOUHDJJ3IrqS02
l57/NPSjNU1Iwd8iM8VOjycPo9F64wxdaILWL0k3Q7kyaeN4Po5rgPYqm49dzxYBQPk1JIkrQ2tA
SCY7OhbPsqlDZ34QK6/jAOs41lANul9aPRl80/IZrKxcuTGwFc3oTDQDHJk0kwMfZfp0ZMb4FkPT
Ct91J8Jn9SFIyDcLld4W8b/nK4KGuXogAMqhAkAwM+EXSVlGWzghSz/TLeKycxBZxiE5vK4A3ZQF
NVu1roT8sfH1RV+INI9k1cAX2gG/rf7Pdj/Z0G+6FL7fY8AIpSfLiAWDrjp8lezrUDps48v4F7Ct
G1s8JLbrGjCFJRq5cRjfXsx/GW5ZwJL3LGZ9txMwSFa9wg1p6NdgVwqDjc0G0INe2CN12ch9qgzf
kzJjDcA3KcY6lr2yaFBHghE5MmBtVZRm7KOvpDlEoBvHoBOax5xrsQ3F8BNs8Dkup4DPND4STW57
AqM62YV0kykH+z6hnAU/U73PFRZ2lszn45PCvLDgX/7rtOw1KlFU140i73YWfWnk673zvIVRxdcx
xHxVv0CfRlrecokAysJyFbiqqdP/Xa34pPcrUCsU/bdjySrCofu6+8SXxJCpm1xfKuuw7g8XTjRb
TWrJmA9efqN0P79dbmOD3qJm2nFOtaU4aO5O/uY80JKe8bxTsb7fwL7Hvr9519fT1K/RkAJCRPHm
M/gpzQdtQrUpdK4fQ2k1XoIBjTET7XRQR+5csGaD1ZH7da0arOV3HHKiA31pYBX+NMg1FcCUdifp
TqBdTtOz9DtpsVRNw8DHaCb10mB8lQJ+C9usbIw/G8Qwuv5YZ6mSRrfdjxPl3by5prKyKBMx1mOH
mVKFtaJi
`pragma protect end_protected

