`timescale 1ns / 1ns
`define SYNTH
//////////////////////////////////////////////////////////////////////////////////
// Company: 浪潮信息
// Engineer: 邓子为
//////////////////////////////////////////////////////////////////////////////////

module top #(
  parameter SIZE_LOOP = 128  //计算的平面数量
  ) (
`ifdef SYNTH
  input         init_clk,      //初始化时钟
  input         sys_clk_clk_p, //PCIe时钟
  input         sys_clk_clk_n,
  input         sys_rstn,      //PCIe复位
  input  [15:0] pcie_mgt_rxn,  //PCIe引脚
  input  [15:0] pcie_mgt_rxp,
  output [15:0] pcie_mgt_txn,
  output [15:0] pcie_mgt_txp
`else
  input         sclk,  
  input         xdma_rstn, 
  input  [31:0] gpio
`endif
);

localparam LENGTH      = 128; //FFT的点数
localparam FFT_NUM     = 8;  //FFT核数量
localparam DWIDTH_FFT  = 32; //FFT数据实部和虚部位宽，BIT
localparam DWIDTH_BRAM = 64; //本地内存的数据位宽，BIT
localparam AWIDTH_BRAM = 14; //本地内存的地址位宽
localparam AWIDTH_HBM  = 32; //全局内存的地址位宽
localparam DWIDTH_HBM  = 32; //全局内存的数据位宽，BYTE
localparam DWIDTH_LOAD = 64; //LOAD模块读数据位宽，BYTE
localparam NUM_GROUP   = 16;  //分组数量
localparam SIZE_GROUP  = LENGTH/NUM_GROUP;

/**************************** XDMA系统 ****************************/
wire    [NUM_GROUP-1:0] s_axi_awready;
wire    [NUM_GROUP-1:0] s_axi_awvalid;
wire   [AWIDTH_HBM-1:0] s_axi_awaddr  [NUM_GROUP-1:0];
wire              [1:0] s_axi_awburst [NUM_GROUP-1:0];
wire              [3:0] s_axi_awcache [NUM_GROUP-1:0];
wire              [7:0] s_axi_awlen   [NUM_GROUP-1:0];
wire              [2:0] s_axi_awsize  [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] s_axi_wready;
wire    [NUM_GROUP-1:0] s_axi_wvalid;
wire [DWIDTH_HBM*8-1:0] s_axi_wdata   [NUM_GROUP-1:0];
wire   [DWIDTH_HBM-1:0] s_axi_wstrb   [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] s_axi_wlast;
wire    [NUM_GROUP-1:0] s_axi_bready;
wire    [NUM_GROUP-1:0] s_axi_bvalid;
wire              [1:0] s_axi_bresp   [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] s_axi_arready;
wire    [NUM_GROUP-1:0] s_axi_arvalid;
wire   [AWIDTH_HBM-1:0] s_axi_araddr  [NUM_GROUP-1:0];
wire              [1:0] s_axi_arburst [NUM_GROUP-1:0];
wire              [3:0] s_axi_arcache [NUM_GROUP-1:0];
wire              [7:0] s_axi_arlen   [NUM_GROUP-1:0];
wire              [2:0] s_axi_arsize  [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] s_axi_rready;
wire    [NUM_GROUP-1:0] s_axi_rvalid;
wire [DWIDTH_HBM*8-1:0] s_axi_rdata   [NUM_GROUP-1:0];
wire    [NUM_GROUP-1:0] s_axi_rlast;
wire              [1:0] s_axi_rresp   [NUM_GROUP-1:0];

wire     [NUM_GROUP-1:0] m_axi_awready;
wire     [NUM_GROUP-1:0] m_axi_awvalid;
wire    [AWIDTH_HBM-1:0] m_axi_awaddr  [NUM_GROUP-1:0];
wire               [1:0] m_axi_awburst [NUM_GROUP-1:0];
wire               [3:0] m_axi_awcache [NUM_GROUP-1:0];
wire               [7:0] m_axi_awlen   [NUM_GROUP-1:0];
wire               [2:0] m_axi_awsize  [NUM_GROUP-1:0];
wire     [NUM_GROUP-1:0] m_axi_wready;
wire     [NUM_GROUP-1:0] m_axi_wvalid;
wire [DWIDTH_LOAD*8-1:0] m_axi_wdata   [NUM_GROUP-1:0];
wire   [DWIDTH_LOAD-1:0] m_axi_wstrb   [NUM_GROUP-1:0];
wire     [NUM_GROUP-1:0] m_axi_wlast;
wire     [NUM_GROUP-1:0] m_axi_bready;
wire     [NUM_GROUP-1:0] m_axi_bvalid;
wire               [1:0] m_axi_bresp   [NUM_GROUP-1:0];
wire     [NUM_GROUP-1:0] m_axi_arready;
wire     [NUM_GROUP-1:0] m_axi_arvalid;
wire    [AWIDTH_HBM-1:0] m_axi_araddr  [NUM_GROUP-1:0];
wire               [1:0] m_axi_arburst [NUM_GROUP-1:0];
wire               [3:0] m_axi_arcache [NUM_GROUP-1:0];
wire               [7:0] m_axi_arlen   [NUM_GROUP-1:0];
wire               [2:0] m_axi_arsize  [NUM_GROUP-1:0];
wire     [NUM_GROUP-1:0] m_axi_rready;
wire     [NUM_GROUP-1:0] m_axi_rvalid;
wire [DWIDTH_LOAD*8-1:0] m_axi_rdata   [NUM_GROUP-1:0];
wire     [NUM_GROUP-1:0] m_axi_rlast;
wire               [1:0] m_axi_rresp   [NUM_GROUP-1:0];

`ifdef SYNTH
wire [31:0] gpio;
xdma_wrapper xdma_wrapper_i(
  .hbm_refclk     (init_clk),
  .pcie_mgt_rxn   (pcie_mgt_rxn),
  .pcie_mgt_rxp   (pcie_mgt_rxp),
  .pcie_mgt_txn   (pcie_mgt_txn),
  .pcie_mgt_txp   (pcie_mgt_txp),
  .sys_clk_clk_n  (sys_clk_clk_n),
  .sys_clk_clk_p  (sys_clk_clk_p),
  .sys_rstn       (sys_rstn),
  .xdma_aclk      (sclk),
  .xdma_rstn      (xdma_rstn),
  .hbm_aclk       (hbm_aclk),
  .gpio           (gpio), 
  .msi_enable     (msi_enable),
  .irq_req        (irq_req),

  .cu_axi0_awready (s_axi_awready[0]),
  .cu_axi0_awvalid (s_axi_awvalid[0]),
  .cu_axi0_awaddr  (s_axi_awaddr [0]),
  .cu_axi0_wready  (s_axi_wready [0]),
  .cu_axi0_wvalid  (s_axi_wvalid [0]),
  .cu_axi0_wdata   (s_axi_wdata  [0]),
  .cu_axi0_wstrb   (s_axi_wstrb  [0]),
  .cu_axi0_wlast   (s_axi_wlast  [0]),
  .cu_axi0_bready  (s_axi_bready [0]),
  .cu_axi0_bvalid  (s_axi_bvalid [0]),
  .cu_axi0_bresp   (s_axi_bresp  [0]),
  .cu_axi0_awburst (s_axi_awburst[0]),
  .cu_axi0_awcache (s_axi_awcache[0]),
  .cu_axi0_awlen   (s_axi_awlen  [0]),
  .cu_axi0_awsize  (s_axi_awsize [0]),
  .cu_axi0_arready (s_axi_arready[0]),
  .cu_axi0_arvalid (s_axi_arvalid[0]),
  .cu_axi0_araddr  (s_axi_araddr [0]),
  .cu_axi0_rready  (s_axi_rready [0]),
  .cu_axi0_rvalid  (s_axi_rvalid [0]),
  .cu_axi0_rdata   (s_axi_rdata  [0]),
  .cu_axi0_rlast   (s_axi_rlast  [0]),
  .cu_axi0_rresp   (s_axi_rresp  [0]),
  .cu_axi0_arburst (s_axi_arburst[0]),
  .cu_axi0_arcache (s_axi_arcache[0]),
  .cu_axi0_arlen   (s_axi_arlen  [0]),
  .cu_axi0_arsize  (s_axi_arsize [0]),
  .cu_axi0_awprot  (),
  .cu_axi0_awlock  (),
  .cu_axi0_awqos   (),
  .cu_axi0_awregion(),
  .cu_axi0_arprot  (),
  .cu_axi0_arlock  (),
  .cu_axi0_arqos   (),
  .cu_axi0_arregion(),

  .cu_axi1_awready (s_axi_awready[1]),
  .cu_axi1_awvalid (s_axi_awvalid[1]),
  .cu_axi1_awaddr  (s_axi_awaddr [1]),
  .cu_axi1_wready  (s_axi_wready [1]),
  .cu_axi1_wvalid  (s_axi_wvalid [1]),
  .cu_axi1_wdata   (s_axi_wdata  [1]),
  .cu_axi1_wstrb   (s_axi_wstrb  [1]),
  .cu_axi1_wlast   (s_axi_wlast  [1]),
  .cu_axi1_bready  (s_axi_bready [1]),
  .cu_axi1_bvalid  (s_axi_bvalid [1]),
  .cu_axi1_bresp   (s_axi_bresp  [1]),
  .cu_axi1_awburst (s_axi_awburst[1]),
  .cu_axi1_awcache (s_axi_awcache[1]),
  .cu_axi1_awlen   (s_axi_awlen  [1]),
  .cu_axi1_awsize  (s_axi_awsize [1]),
  .cu_axi1_arready (s_axi_arready[1]),
  .cu_axi1_arvalid (s_axi_arvalid[1]),
  .cu_axi1_araddr  (s_axi_araddr [1]),
  .cu_axi1_rready  (s_axi_rready [1]),
  .cu_axi1_rvalid  (s_axi_rvalid [1]),
  .cu_axi1_rdata   (s_axi_rdata  [1]),
  .cu_axi1_rlast   (s_axi_rlast  [1]),
  .cu_axi1_rresp   (s_axi_rresp  [1]),
  .cu_axi1_arburst (s_axi_arburst[1]),
  .cu_axi1_arcache (s_axi_arcache[1]),
  .cu_axi1_arlen   (s_axi_arlen  [1]),
  .cu_axi1_arsize  (s_axi_arsize [1]),
  .cu_axi1_awprot  (),
  .cu_axi1_awlock  (),
  .cu_axi1_awqos   (),
  .cu_axi1_awregion(),
  .cu_axi1_arprot  (),
  .cu_axi1_arlock  (),
  .cu_axi1_arqos   (),
  .cu_axi1_arregion(),

  .cu_axi2_awready (s_axi_awready[2]),
  .cu_axi2_awvalid (s_axi_awvalid[2]),
  .cu_axi2_awaddr  (s_axi_awaddr [2]),
  .cu_axi2_wready  (s_axi_wready [2]),
  .cu_axi2_wvalid  (s_axi_wvalid [2]),
  .cu_axi2_wdata   (s_axi_wdata  [2]),
  .cu_axi2_wstrb   (s_axi_wstrb  [2]),
  .cu_axi2_wlast   (s_axi_wlast  [2]),
  .cu_axi2_bready  (s_axi_bready [2]),
  .cu_axi2_bvalid  (s_axi_bvalid [2]),
  .cu_axi2_bresp   (s_axi_bresp  [2]),
  .cu_axi2_awburst (s_axi_awburst[2]),
  .cu_axi2_awcache (s_axi_awcache[2]),
  .cu_axi2_awlen   (s_axi_awlen  [2]),
  .cu_axi2_awsize  (s_axi_awsize [2]),
  .cu_axi2_arready (s_axi_arready[2]),
  .cu_axi2_arvalid (s_axi_arvalid[2]),
  .cu_axi2_araddr  (s_axi_araddr [2]),
  .cu_axi2_rready  (s_axi_rready [2]),
  .cu_axi2_rvalid  (s_axi_rvalid [2]),
  .cu_axi2_rdata   (s_axi_rdata  [2]),
  .cu_axi2_rlast   (s_axi_rlast  [2]),
  .cu_axi2_rresp   (s_axi_rresp  [2]),
  .cu_axi2_arburst (s_axi_arburst[2]),
  .cu_axi2_arcache (s_axi_arcache[2]),
  .cu_axi2_arlen   (s_axi_arlen  [2]),
  .cu_axi2_arsize  (s_axi_arsize [2]),
  .cu_axi2_awprot  (),
  .cu_axi2_awlock  (),
  .cu_axi2_awqos   (),
  .cu_axi2_awregion(),
  .cu_axi2_arprot  (),
  .cu_axi2_arlock  (),
  .cu_axi2_arqos   (),
  .cu_axi2_arregion(),

  .cu_axi3_awready (s_axi_awready[3]),
  .cu_axi3_awvalid (s_axi_awvalid[3]),
  .cu_axi3_awaddr  (s_axi_awaddr [3]),
  .cu_axi3_wready  (s_axi_wready [3]),
  .cu_axi3_wvalid  (s_axi_wvalid [3]),
  .cu_axi3_wdata   (s_axi_wdata  [3]),
  .cu_axi3_wstrb   (s_axi_wstrb  [3]),
  .cu_axi3_wlast   (s_axi_wlast  [3]),
  .cu_axi3_bready  (s_axi_bready [3]),
  .cu_axi3_bvalid  (s_axi_bvalid [3]),
  .cu_axi3_bresp   (s_axi_bresp  [3]),
  .cu_axi3_awburst (s_axi_awburst[3]),
  .cu_axi3_awcache (s_axi_awcache[3]),
  .cu_axi3_awlen   (s_axi_awlen  [3]),
  .cu_axi3_awsize  (s_axi_awsize [3]),
  .cu_axi3_arready (s_axi_arready[3]),
  .cu_axi3_arvalid (s_axi_arvalid[3]),
  .cu_axi3_araddr  (s_axi_araddr [3]),
  .cu_axi3_rready  (s_axi_rready [3]),
  .cu_axi3_rvalid  (s_axi_rvalid [3]),
  .cu_axi3_rdata   (s_axi_rdata  [3]),
  .cu_axi3_rlast   (s_axi_rlast  [3]),
  .cu_axi3_rresp   (s_axi_rresp  [3]),
  .cu_axi3_arburst (s_axi_arburst[3]),
  .cu_axi3_arcache (s_axi_arcache[3]),
  .cu_axi3_arlen   (s_axi_arlen  [3]),
  .cu_axi3_arsize  (s_axi_arsize [3]),
  .cu_axi3_awprot  (),
  .cu_axi3_awlock  (),
  .cu_axi3_awqos   (),
  .cu_axi3_awregion(),
  .cu_axi3_arprot  (),
  .cu_axi3_arlock  (),
  .cu_axi3_arqos   (),
  .cu_axi3_arregion(),

  .cu_axi4_awready (s_axi_awready[4]),
  .cu_axi4_awvalid (s_axi_awvalid[4]),
  .cu_axi4_awaddr  (s_axi_awaddr [4]),
  .cu_axi4_wready  (s_axi_wready [4]),
  .cu_axi4_wvalid  (s_axi_wvalid [4]),
  .cu_axi4_wdata   (s_axi_wdata  [4]),
  .cu_axi4_wstrb   (s_axi_wstrb  [4]),
  .cu_axi4_wlast   (s_axi_wlast  [4]),
  .cu_axi4_bready  (s_axi_bready [4]),
  .cu_axi4_bvalid  (s_axi_bvalid [4]),
  .cu_axi4_bresp   (s_axi_bresp  [4]),
  .cu_axi4_awburst (s_axi_awburst[4]),
  .cu_axi4_awcache (s_axi_awcache[4]),
  .cu_axi4_awlen   (s_axi_awlen  [4]),
  .cu_axi4_awsize  (s_axi_awsize [4]),
  .cu_axi4_arready (s_axi_arready[4]),
  .cu_axi4_arvalid (s_axi_arvalid[4]),
  .cu_axi4_araddr  (s_axi_araddr [4]),
  .cu_axi4_rready  (s_axi_rready [4]),
  .cu_axi4_rvalid  (s_axi_rvalid [4]),
  .cu_axi4_rdata   (s_axi_rdata  [4]),
  .cu_axi4_rlast   (s_axi_rlast  [4]),
  .cu_axi4_rresp   (s_axi_rresp  [4]),
  .cu_axi4_arburst (s_axi_arburst[4]),
  .cu_axi4_arcache (s_axi_arcache[4]),
  .cu_axi4_arlen   (s_axi_arlen  [4]),
  .cu_axi4_arsize  (s_axi_arsize [4]),
  .cu_axi4_awprot  (),
  .cu_axi4_awlock  (),
  .cu_axi4_awqos   (),
  .cu_axi4_awregion(),
  .cu_axi4_arprot  (),
  .cu_axi4_arlock  (),
  .cu_axi4_arqos   (),
  .cu_axi4_arregion(),

  .cu_axi5_awready (s_axi_awready[5]),
  .cu_axi5_awvalid (s_axi_awvalid[5]),
  .cu_axi5_awaddr  (s_axi_awaddr [5]),
  .cu_axi5_wready  (s_axi_wready [5]),
  .cu_axi5_wvalid  (s_axi_wvalid [5]),
  .cu_axi5_wdata   (s_axi_wdata  [5]),
  .cu_axi5_wstrb   (s_axi_wstrb  [5]),
  .cu_axi5_wlast   (s_axi_wlast  [5]),
  .cu_axi5_bready  (s_axi_bready [5]),
  .cu_axi5_bvalid  (s_axi_bvalid [5]),
  .cu_axi5_bresp   (s_axi_bresp  [5]),
  .cu_axi5_awburst (s_axi_awburst[5]),
  .cu_axi5_awcache (s_axi_awcache[5]),
  .cu_axi5_awlen   (s_axi_awlen  [5]),
  .cu_axi5_awsize  (s_axi_awsize [5]),
  .cu_axi5_arready (s_axi_arready[5]),
  .cu_axi5_arvalid (s_axi_arvalid[5]),
  .cu_axi5_araddr  (s_axi_araddr [5]),
  .cu_axi5_rready  (s_axi_rready [5]),
  .cu_axi5_rvalid  (s_axi_rvalid [5]),
  .cu_axi5_rdata   (s_axi_rdata  [5]),
  .cu_axi5_rlast   (s_axi_rlast  [5]),
  .cu_axi5_rresp   (s_axi_rresp  [5]),
  .cu_axi5_arburst (s_axi_arburst[5]),
  .cu_axi5_arcache (s_axi_arcache[5]),
  .cu_axi5_arlen   (s_axi_arlen  [5]),
  .cu_axi5_arsize  (s_axi_arsize [5]),
  .cu_axi5_awprot  (),
  .cu_axi5_awlock  (),
  .cu_axi5_awqos   (),
  .cu_axi5_awregion(),
  .cu_axi5_arprot  (),
  .cu_axi5_arlock  (),
  .cu_axi5_arqos   (),
  .cu_axi5_arregion(),

  .cu_axi6_awready (s_axi_awready[6]),
  .cu_axi6_awvalid (s_axi_awvalid[6]),
  .cu_axi6_awaddr  (s_axi_awaddr [6]),
  .cu_axi6_wready  (s_axi_wready [6]),
  .cu_axi6_wvalid  (s_axi_wvalid [6]),
  .cu_axi6_wdata   (s_axi_wdata  [6]),
  .cu_axi6_wstrb   (s_axi_wstrb  [6]),
  .cu_axi6_wlast   (s_axi_wlast  [6]),
  .cu_axi6_bready  (s_axi_bready [6]),
  .cu_axi6_bvalid  (s_axi_bvalid [6]),
  .cu_axi6_bresp   (s_axi_bresp  [6]),
  .cu_axi6_awburst (s_axi_awburst[6]),
  .cu_axi6_awcache (s_axi_awcache[6]),
  .cu_axi6_awlen   (s_axi_awlen  [6]),
  .cu_axi6_awsize  (s_axi_awsize [6]),
  .cu_axi6_arready (s_axi_arready[6]),
  .cu_axi6_arvalid (s_axi_arvalid[6]),
  .cu_axi6_araddr  (s_axi_araddr [6]),
  .cu_axi6_rready  (s_axi_rready [6]),
  .cu_axi6_rvalid  (s_axi_rvalid [6]),
  .cu_axi6_rdata   (s_axi_rdata  [6]),
  .cu_axi6_rlast   (s_axi_rlast  [6]),
  .cu_axi6_rresp   (s_axi_rresp  [6]),
  .cu_axi6_arburst (s_axi_arburst[6]),
  .cu_axi6_arcache (s_axi_arcache[6]),
  .cu_axi6_arlen   (s_axi_arlen  [6]),
  .cu_axi6_arsize  (s_axi_arsize [6]),
  .cu_axi6_awprot  (),
  .cu_axi6_awlock  (),
  .cu_axi6_awqos   (),
  .cu_axi6_awregion(),
  .cu_axi6_arprot  (),
  .cu_axi6_arlock  (),
  .cu_axi6_arqos   (),
  .cu_axi6_arregion(),

  .cu_axi7_awready (s_axi_awready[7]),
  .cu_axi7_awvalid (s_axi_awvalid[7]),
  .cu_axi7_awaddr  (s_axi_awaddr [7]),
  .cu_axi7_wready  (s_axi_wready [7]),
  .cu_axi7_wvalid  (s_axi_wvalid [7]),
  .cu_axi7_wdata   (s_axi_wdata  [7]),
  .cu_axi7_wstrb   (s_axi_wstrb  [7]),
  .cu_axi7_wlast   (s_axi_wlast  [7]),
  .cu_axi7_bready  (s_axi_bready [7]),
  .cu_axi7_bvalid  (s_axi_bvalid [7]),
  .cu_axi7_bresp   (s_axi_bresp  [7]),
  .cu_axi7_awburst (s_axi_awburst[7]),
  .cu_axi7_awcache (s_axi_awcache[7]),
  .cu_axi7_awlen   (s_axi_awlen  [7]),
  .cu_axi7_awsize  (s_axi_awsize [7]),
  .cu_axi7_arready (s_axi_arready[7]),
  .cu_axi7_arvalid (s_axi_arvalid[7]),
  .cu_axi7_araddr  (s_axi_araddr [7]),
  .cu_axi7_rready  (s_axi_rready [7]),
  .cu_axi7_rvalid  (s_axi_rvalid [7]),
  .cu_axi7_rdata   (s_axi_rdata  [7]),
  .cu_axi7_rlast   (s_axi_rlast  [7]),
  .cu_axi7_rresp   (s_axi_rresp  [7]),
  .cu_axi7_arburst (s_axi_arburst[7]),
  .cu_axi7_arcache (s_axi_arcache[7]),
  .cu_axi7_arlen   (s_axi_arlen  [7]),
  .cu_axi7_arsize  (s_axi_arsize [7]),
  .cu_axi7_awprot  (),
  .cu_axi7_awlock  (),
  .cu_axi7_awqos   (),
  .cu_axi7_awregion(),
  .cu_axi7_arprot  (),
  .cu_axi7_arlock  (),
  .cu_axi7_arqos   (),
  .cu_axi7_arregion(),

  .cu_axi8_awready (s_axi_awready[8]),
  .cu_axi8_awvalid (s_axi_awvalid[8]),
  .cu_axi8_awaddr  (s_axi_awaddr [8]),
  .cu_axi8_wready  (s_axi_wready [8]),
  .cu_axi8_wvalid  (s_axi_wvalid [8]),
  .cu_axi8_wdata   (s_axi_wdata  [8]),
  .cu_axi8_wstrb   (s_axi_wstrb  [8]),
  .cu_axi8_wlast   (s_axi_wlast  [8]),
  .cu_axi8_bready  (s_axi_bready [8]),
  .cu_axi8_bvalid  (s_axi_bvalid [8]),
  .cu_axi8_bresp   (s_axi_bresp  [8]),
  .cu_axi8_awburst (s_axi_awburst[8]),
  .cu_axi8_awcache (s_axi_awcache[8]),
  .cu_axi8_awlen   (s_axi_awlen  [8]),
  .cu_axi8_awsize  (s_axi_awsize [8]),
  .cu_axi8_arready (s_axi_arready[8]),
  .cu_axi8_arvalid (s_axi_arvalid[8]),
  .cu_axi8_araddr  (s_axi_araddr [8]),
  .cu_axi8_rready  (s_axi_rready [8]),
  .cu_axi8_rvalid  (s_axi_rvalid [8]),
  .cu_axi8_rdata   (s_axi_rdata  [8]),
  .cu_axi8_rlast   (s_axi_rlast  [8]),
  .cu_axi8_rresp   (s_axi_rresp  [8]),
  .cu_axi8_arburst (s_axi_arburst[8]),
  .cu_axi8_arcache (s_axi_arcache[8]),
  .cu_axi8_arlen   (s_axi_arlen  [8]),
  .cu_axi8_arsize  (s_axi_arsize [8]),
  .cu_axi8_awprot  (),
  .cu_axi8_awlock  (),
  .cu_axi8_awqos   (),
  .cu_axi8_awregion(),
  .cu_axi8_arprot  (),
  .cu_axi8_arlock  (),
  .cu_axi8_arqos   (),
  .cu_axi8_arregion(),

  .cu_axi9_awready (s_axi_awready[9]),
  .cu_axi9_awvalid (s_axi_awvalid[9]),
  .cu_axi9_awaddr  (s_axi_awaddr [9]),
  .cu_axi9_wready  (s_axi_wready [9]),
  .cu_axi9_wvalid  (s_axi_wvalid [9]),
  .cu_axi9_wdata   (s_axi_wdata  [9]),
  .cu_axi9_wstrb   (s_axi_wstrb  [9]),
  .cu_axi9_wlast   (s_axi_wlast  [9]),
  .cu_axi9_bready  (s_axi_bready [9]),
  .cu_axi9_bvalid  (s_axi_bvalid [9]),
  .cu_axi9_bresp   (s_axi_bresp  [9]),
  .cu_axi9_awburst (s_axi_awburst[9]),
  .cu_axi9_awcache (s_axi_awcache[9]),
  .cu_axi9_awlen   (s_axi_awlen  [9]),
  .cu_axi9_awsize  (s_axi_awsize [9]),
  .cu_axi9_arready (s_axi_arready[9]),
  .cu_axi9_arvalid (s_axi_arvalid[9]),
  .cu_axi9_araddr  (s_axi_araddr [9]),
  .cu_axi9_rready  (s_axi_rready [9]),
  .cu_axi9_rvalid  (s_axi_rvalid [9]),
  .cu_axi9_rdata   (s_axi_rdata  [9]),
  .cu_axi9_rlast   (s_axi_rlast  [9]),
  .cu_axi9_rresp   (s_axi_rresp  [9]),
  .cu_axi9_arburst (s_axi_arburst[9]),
  .cu_axi9_arcache (s_axi_arcache[9]),
  .cu_axi9_arlen   (s_axi_arlen  [9]),
  .cu_axi9_arsize  (s_axi_arsize [9]),
  .cu_axi9_awprot  (),
  .cu_axi9_awlock  (),
  .cu_axi9_awqos   (),
  .cu_axi9_awregion(),
  .cu_axi9_arprot  (),
  .cu_axi9_arlock  (),
  .cu_axi9_arqos   (),
  .cu_axi9_arregion(),

  .cu_axi10_awready (s_axi_awready[10]),
  .cu_axi10_awvalid (s_axi_awvalid[10]),
  .cu_axi10_awaddr  (s_axi_awaddr [10]),
  .cu_axi10_wready  (s_axi_wready [10]),
  .cu_axi10_wvalid  (s_axi_wvalid [10]),
  .cu_axi10_wdata   (s_axi_wdata  [10]),
  .cu_axi10_wstrb   (s_axi_wstrb  [10]),
  .cu_axi10_wlast   (s_axi_wlast  [10]),
  .cu_axi10_bready  (s_axi_bready [10]),
  .cu_axi10_bvalid  (s_axi_bvalid [10]),
  .cu_axi10_bresp   (s_axi_bresp  [10]),
  .cu_axi10_awburst (s_axi_awburst[10]),
  .cu_axi10_awcache (s_axi_awcache[10]),
  .cu_axi10_awlen   (s_axi_awlen  [10]),
  .cu_axi10_awsize  (s_axi_awsize [10]),
  .cu_axi10_arready (s_axi_arready[10]),
  .cu_axi10_arvalid (s_axi_arvalid[10]),
  .cu_axi10_araddr  (s_axi_araddr [10]),
  .cu_axi10_rready  (s_axi_rready [10]),
  .cu_axi10_rvalid  (s_axi_rvalid [10]),
  .cu_axi10_rdata   (s_axi_rdata  [10]),
  .cu_axi10_rlast   (s_axi_rlast  [10]),
  .cu_axi10_rresp   (s_axi_rresp  [10]),
  .cu_axi10_arburst (s_axi_arburst[10]),
  .cu_axi10_arcache (s_axi_arcache[10]),
  .cu_axi10_arlen   (s_axi_arlen  [10]),
  .cu_axi10_arsize  (s_axi_arsize [10]),
  .cu_axi10_awprot  (),
  .cu_axi10_awlock  (),
  .cu_axi10_awqos   (),
  .cu_axi10_awregion(),
  .cu_axi10_arprot  (),
  .cu_axi10_arlock  (),
  .cu_axi10_arqos   (),
  .cu_axi10_arregion(),

  .cu_axi11_awready (s_axi_awready[11]),
  .cu_axi11_awvalid (s_axi_awvalid[11]),
  .cu_axi11_awaddr  (s_axi_awaddr [11]),
  .cu_axi11_wready  (s_axi_wready [11]),
  .cu_axi11_wvalid  (s_axi_wvalid [11]),
  .cu_axi11_wdata   (s_axi_wdata  [11]),
  .cu_axi11_wstrb   (s_axi_wstrb  [11]),
  .cu_axi11_wlast   (s_axi_wlast  [11]),
  .cu_axi11_bready  (s_axi_bready [11]),
  .cu_axi11_bvalid  (s_axi_bvalid [11]),
  .cu_axi11_bresp   (s_axi_bresp  [11]),
  .cu_axi11_awburst (s_axi_awburst[11]),
  .cu_axi11_awcache (s_axi_awcache[11]),
  .cu_axi11_awlen   (s_axi_awlen  [11]),
  .cu_axi11_awsize  (s_axi_awsize [11]),
  .cu_axi11_arready (s_axi_arready[11]),
  .cu_axi11_arvalid (s_axi_arvalid[11]),
  .cu_axi11_araddr  (s_axi_araddr [11]),
  .cu_axi11_rready  (s_axi_rready [11]),
  .cu_axi11_rvalid  (s_axi_rvalid [11]),
  .cu_axi11_rdata   (s_axi_rdata  [11]),
  .cu_axi11_rlast   (s_axi_rlast  [11]),
  .cu_axi11_rresp   (s_axi_rresp  [11]),
  .cu_axi11_arburst (s_axi_arburst[11]),
  .cu_axi11_arcache (s_axi_arcache[11]),
  .cu_axi11_arlen   (s_axi_arlen  [11]),
  .cu_axi11_arsize  (s_axi_arsize [11]),
  .cu_axi11_awprot  (),
  .cu_axi11_awlock  (),
  .cu_axi11_awqos   (),
  .cu_axi11_awregion(),
  .cu_axi11_arprot  (),
  .cu_axi11_arlock  (),
  .cu_axi11_arqos   (),
  .cu_axi11_arregion(),

  .cu_axi12_awready (s_axi_awready[12]),
  .cu_axi12_awvalid (s_axi_awvalid[12]),
  .cu_axi12_awaddr  (s_axi_awaddr [12]),
  .cu_axi12_wready  (s_axi_wready [12]),
  .cu_axi12_wvalid  (s_axi_wvalid [12]),
  .cu_axi12_wdata   (s_axi_wdata  [12]),
  .cu_axi12_wstrb   (s_axi_wstrb  [12]),
  .cu_axi12_wlast   (s_axi_wlast  [12]),
  .cu_axi12_bready  (s_axi_bready [12]),
  .cu_axi12_bvalid  (s_axi_bvalid [12]),
  .cu_axi12_bresp   (s_axi_bresp  [12]),
  .cu_axi12_awburst (s_axi_awburst[12]),
  .cu_axi12_awcache (s_axi_awcache[12]),
  .cu_axi12_awlen   (s_axi_awlen  [12]),
  .cu_axi12_awsize  (s_axi_awsize [12]),
  .cu_axi12_arready (s_axi_arready[12]),
  .cu_axi12_arvalid (s_axi_arvalid[12]),
  .cu_axi12_araddr  (s_axi_araddr [12]),
  .cu_axi12_rready  (s_axi_rready [12]),
  .cu_axi12_rvalid  (s_axi_rvalid [12]),
  .cu_axi12_rdata   (s_axi_rdata  [12]),
  .cu_axi12_rlast   (s_axi_rlast  [12]),
  .cu_axi12_rresp   (s_axi_rresp  [12]),
  .cu_axi12_arburst (s_axi_arburst[12]),
  .cu_axi12_arcache (s_axi_arcache[12]),
  .cu_axi12_arlen   (s_axi_arlen  [12]),
  .cu_axi12_arsize  (s_axi_arsize [12]),
  .cu_axi12_awprot  (),
  .cu_axi12_awlock  (),
  .cu_axi12_awqos   (),
  .cu_axi12_awregion(),
  .cu_axi12_arprot  (),
  .cu_axi12_arlock  (),
  .cu_axi12_arqos   (),
  .cu_axi12_arregion(),

  .cu_axi13_awready (s_axi_awready[13]),
  .cu_axi13_awvalid (s_axi_awvalid[13]),
  .cu_axi13_awaddr  (s_axi_awaddr [13]),
  .cu_axi13_wready  (s_axi_wready [13]),
  .cu_axi13_wvalid  (s_axi_wvalid [13]),
  .cu_axi13_wdata   (s_axi_wdata  [13]),
  .cu_axi13_wstrb   (s_axi_wstrb  [13]),
  .cu_axi13_wlast   (s_axi_wlast  [13]),
  .cu_axi13_bready  (s_axi_bready [13]),
  .cu_axi13_bvalid  (s_axi_bvalid [13]),
  .cu_axi13_bresp   (s_axi_bresp  [13]),
  .cu_axi13_awburst (s_axi_awburst[13]),
  .cu_axi13_awcache (s_axi_awcache[13]),
  .cu_axi13_awlen   (s_axi_awlen  [13]),
  .cu_axi13_awsize  (s_axi_awsize [13]),
  .cu_axi13_arready (s_axi_arready[13]),
  .cu_axi13_arvalid (s_axi_arvalid[13]),
  .cu_axi13_araddr  (s_axi_araddr [13]),
  .cu_axi13_rready  (s_axi_rready [13]),
  .cu_axi13_rvalid  (s_axi_rvalid [13]),
  .cu_axi13_rdata   (s_axi_rdata  [13]),
  .cu_axi13_rlast   (s_axi_rlast  [13]),
  .cu_axi13_rresp   (s_axi_rresp  [13]),
  .cu_axi13_arburst (s_axi_arburst[13]),
  .cu_axi13_arcache (s_axi_arcache[13]),
  .cu_axi13_arlen   (s_axi_arlen  [13]),
  .cu_axi13_arsize  (s_axi_arsize [13]),
  .cu_axi13_awprot  (),
  .cu_axi13_awlock  (),
  .cu_axi13_awqos   (),
  .cu_axi13_awregion(),
  .cu_axi13_arprot  (),
  .cu_axi13_arlock  (),
  .cu_axi13_arqos   (),
  .cu_axi13_arregion(),

  .cu_axi14_awready (s_axi_awready[14]),
  .cu_axi14_awvalid (s_axi_awvalid[14]),
  .cu_axi14_awaddr  (s_axi_awaddr [14]),
  .cu_axi14_wready  (s_axi_wready [14]),
  .cu_axi14_wvalid  (s_axi_wvalid [14]),
  .cu_axi14_wdata   (s_axi_wdata  [14]),
  .cu_axi14_wstrb   (s_axi_wstrb  [14]),
  .cu_axi14_wlast   (s_axi_wlast  [14]),
  .cu_axi14_bready  (s_axi_bready [14]),
  .cu_axi14_bvalid  (s_axi_bvalid [14]),
  .cu_axi14_bresp   (s_axi_bresp  [14]),
  .cu_axi14_awburst (s_axi_awburst[14]),
  .cu_axi14_awcache (s_axi_awcache[14]),
  .cu_axi14_awlen   (s_axi_awlen  [14]),
  .cu_axi14_awsize  (s_axi_awsize [14]),
  .cu_axi14_arready (s_axi_arready[14]),
  .cu_axi14_arvalid (s_axi_arvalid[14]),
  .cu_axi14_araddr  (s_axi_araddr [14]),
  .cu_axi14_rready  (s_axi_rready [14]),
  .cu_axi14_rvalid  (s_axi_rvalid [14]),
  .cu_axi14_rdata   (s_axi_rdata  [14]),
  .cu_axi14_rlast   (s_axi_rlast  [14]),
  .cu_axi14_rresp   (s_axi_rresp  [14]),
  .cu_axi14_arburst (s_axi_arburst[14]),
  .cu_axi14_arcache (s_axi_arcache[14]),
  .cu_axi14_arlen   (s_axi_arlen  [14]),
  .cu_axi14_arsize  (s_axi_arsize [14]),
  .cu_axi14_awprot  (),
  .cu_axi14_awlock  (),
  .cu_axi14_awqos   (),
  .cu_axi14_awregion(),
  .cu_axi14_arprot  (),
  .cu_axi14_arlock  (),
  .cu_axi14_arqos   (),
  .cu_axi14_arregion(),

  .cu_axi15_awready (s_axi_awready[15]),
  .cu_axi15_awvalid (s_axi_awvalid[15]),
  .cu_axi15_awaddr  (s_axi_awaddr [15]),
  .cu_axi15_wready  (s_axi_wready [15]),
  .cu_axi15_wvalid  (s_axi_wvalid [15]),
  .cu_axi15_wdata   (s_axi_wdata  [15]),
  .cu_axi15_wstrb   (s_axi_wstrb  [15]),
  .cu_axi15_wlast   (s_axi_wlast  [15]),
  .cu_axi15_bready  (s_axi_bready [15]),
  .cu_axi15_bvalid  (s_axi_bvalid [15]),
  .cu_axi15_bresp   (s_axi_bresp  [15]),
  .cu_axi15_awburst (s_axi_awburst[15]),
  .cu_axi15_awcache (s_axi_awcache[15]),
  .cu_axi15_awlen   (s_axi_awlen  [15]),
  .cu_axi15_awsize  (s_axi_awsize [15]),
  .cu_axi15_arready (s_axi_arready[15]),
  .cu_axi15_arvalid (s_axi_arvalid[15]),
  .cu_axi15_araddr  (s_axi_araddr [15]),
  .cu_axi15_rready  (s_axi_rready [15]),
  .cu_axi15_rvalid  (s_axi_rvalid [15]),
  .cu_axi15_rdata   (s_axi_rdata  [15]),
  .cu_axi15_rlast   (s_axi_rlast  [15]),
  .cu_axi15_rresp   (s_axi_rresp  [15]),
  .cu_axi15_arburst (s_axi_arburst[15]),
  .cu_axi15_arcache (s_axi_arcache[15]),
  .cu_axi15_arlen   (s_axi_arlen  [15]),
  .cu_axi15_arsize  (s_axi_arsize [15]),
  .cu_axi15_awprot  (),
  .cu_axi15_awlock  (),
  .cu_axi15_awqos   (),
  .cu_axi15_awregion(),
  .cu_axi15_arprot  (),
  .cu_axi15_arlock  (),
  .cu_axi15_arqos   (),
  .cu_axi15_arregion()
);

`else
clkwiz clkwiz_i (
  .clk_in1 (sclk),
  .clk_out1(hbm_aclk)
);

bram_init0 bram0 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[0]),
  .s_axi_awvalid(s_axi_awvalid[0]),
  .s_axi_awaddr (s_axi_awaddr [0]),
  .s_axi_wready (s_axi_wready [0]),
  .s_axi_wvalid (s_axi_wvalid [0]),
  .s_axi_wdata  (s_axi_wdata  [0]),
  .s_axi_wstrb  (s_axi_wstrb  [0]),
  .s_axi_wlast  (s_axi_wlast  [0]),
  .s_axi_bready (s_axi_bready [0]),
  .s_axi_bvalid (s_axi_bvalid [0]),
  .s_axi_bresp  (s_axi_bresp  [0]),
  .s_axi_awlen  (s_axi_awlen  [0]),
  .s_axi_awsize (s_axi_awsize [0]),
  .s_axi_awburst(s_axi_awburst[0]),
  .s_axi_arready(s_axi_arready[0]),
  .s_axi_arvalid(s_axi_arvalid[0]),
  .s_axi_araddr (s_axi_araddr [0]),
  .s_axi_rready (s_axi_rready [0]),
  .s_axi_rvalid (s_axi_rvalid [0]),
  .s_axi_rdata  (s_axi_rdata  [0]),
  .s_axi_rlast  (s_axi_rlast  [0]),
  .s_axi_rresp  (s_axi_rresp  [0]),
  .s_axi_arlen  (s_axi_arlen  [0]),
  .s_axi_arsize (s_axi_arsize [0]),
  .s_axi_arburst(s_axi_arburst[0]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init1 bram1 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[1]),
  .s_axi_awvalid(s_axi_awvalid[1]),
  .s_axi_awaddr (s_axi_awaddr [1]),
  .s_axi_wready (s_axi_wready [1]),
  .s_axi_wvalid (s_axi_wvalid [1]),
  .s_axi_wdata  (s_axi_wdata  [1]),
  .s_axi_wstrb  (s_axi_wstrb  [1]),
  .s_axi_wlast  (s_axi_wlast  [1]),
  .s_axi_bready (s_axi_bready [1]),
  .s_axi_bvalid (s_axi_bvalid [1]),
  .s_axi_bresp  (s_axi_bresp  [1]),
  .s_axi_awlen  (s_axi_awlen  [1]),
  .s_axi_awsize (s_axi_awsize [1]),
  .s_axi_awburst(s_axi_awburst[1]),
  .s_axi_arready(s_axi_arready[1]),
  .s_axi_arvalid(s_axi_arvalid[1]),
  .s_axi_araddr (s_axi_araddr [1]),
  .s_axi_rready (s_axi_rready [1]),
  .s_axi_rvalid (s_axi_rvalid [1]),
  .s_axi_rdata  (s_axi_rdata  [1]),
  .s_axi_rlast  (s_axi_rlast  [1]),
  .s_axi_rresp  (s_axi_rresp  [1]),
  .s_axi_arlen  (s_axi_arlen  [1]),
  .s_axi_arsize (s_axi_arsize [1]),
  .s_axi_arburst(s_axi_arburst[1]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init2 bram2 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[2]),
  .s_axi_awvalid(s_axi_awvalid[2]),
  .s_axi_awaddr (s_axi_awaddr [2]),
  .s_axi_wready (s_axi_wready [2]),
  .s_axi_wvalid (s_axi_wvalid [2]),
  .s_axi_wdata  (s_axi_wdata  [2]),
  .s_axi_wstrb  (s_axi_wstrb  [2]),
  .s_axi_wlast  (s_axi_wlast  [2]),
  .s_axi_bready (s_axi_bready [2]),
  .s_axi_bvalid (s_axi_bvalid [2]),
  .s_axi_bresp  (s_axi_bresp  [2]),
  .s_axi_awlen  (s_axi_awlen  [2]),
  .s_axi_awsize (s_axi_awsize [2]),
  .s_axi_awburst(s_axi_awburst[2]),
  .s_axi_arready(s_axi_arready[2]),
  .s_axi_arvalid(s_axi_arvalid[2]),
  .s_axi_araddr (s_axi_araddr [2]),
  .s_axi_rready (s_axi_rready [2]),
  .s_axi_rvalid (s_axi_rvalid [2]),
  .s_axi_rdata  (s_axi_rdata  [2]),
  .s_axi_rlast  (s_axi_rlast  [2]),
  .s_axi_rresp  (s_axi_rresp  [2]),
  .s_axi_arlen  (s_axi_arlen  [2]),
  .s_axi_arsize (s_axi_arsize [2]),
  .s_axi_arburst(s_axi_arburst[2]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init3 bram3 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[3]),
  .s_axi_awvalid(s_axi_awvalid[3]),
  .s_axi_awaddr (s_axi_awaddr [3]),
  .s_axi_wready (s_axi_wready [3]),
  .s_axi_wvalid (s_axi_wvalid [3]),
  .s_axi_wdata  (s_axi_wdata  [3]),
  .s_axi_wstrb  (s_axi_wstrb  [3]),
  .s_axi_wlast  (s_axi_wlast  [3]),
  .s_axi_bready (s_axi_bready [3]),
  .s_axi_bvalid (s_axi_bvalid [3]),
  .s_axi_bresp  (s_axi_bresp  [3]),
  .s_axi_awlen  (s_axi_awlen  [3]),
  .s_axi_awsize (s_axi_awsize [3]),
  .s_axi_awburst(s_axi_awburst[3]),
  .s_axi_arready(s_axi_arready[3]),
  .s_axi_arvalid(s_axi_arvalid[3]),
  .s_axi_araddr (s_axi_araddr [3]),
  .s_axi_rready (s_axi_rready [3]),
  .s_axi_rvalid (s_axi_rvalid [3]),
  .s_axi_rdata  (s_axi_rdata  [3]),
  .s_axi_rlast  (s_axi_rlast  [3]),
  .s_axi_rresp  (s_axi_rresp  [3]),
  .s_axi_arlen  (s_axi_arlen  [3]),
  .s_axi_arsize (s_axi_arsize [3]),
  .s_axi_arburst(s_axi_arburst[3]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init4 bram4 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[4]),
  .s_axi_awvalid(s_axi_awvalid[4]),
  .s_axi_awaddr (s_axi_awaddr [4]),
  .s_axi_wready (s_axi_wready [4]),
  .s_axi_wvalid (s_axi_wvalid [4]),
  .s_axi_wdata  (s_axi_wdata  [4]),
  .s_axi_wstrb  (s_axi_wstrb  [4]),
  .s_axi_wlast  (s_axi_wlast  [4]),
  .s_axi_bready (s_axi_bready [4]),
  .s_axi_bvalid (s_axi_bvalid [4]),
  .s_axi_bresp  (s_axi_bresp  [4]),
  .s_axi_awlen  (s_axi_awlen  [4]),
  .s_axi_awsize (s_axi_awsize [4]),
  .s_axi_awburst(s_axi_awburst[4]),
  .s_axi_arready(s_axi_arready[4]),
  .s_axi_arvalid(s_axi_arvalid[4]),
  .s_axi_araddr (s_axi_araddr [4]),
  .s_axi_rready (s_axi_rready [4]),
  .s_axi_rvalid (s_axi_rvalid [4]),
  .s_axi_rdata  (s_axi_rdata  [4]),
  .s_axi_rlast  (s_axi_rlast  [4]),
  .s_axi_rresp  (s_axi_rresp  [4]),
  .s_axi_arlen  (s_axi_arlen  [4]),
  .s_axi_arsize (s_axi_arsize [4]),
  .s_axi_arburst(s_axi_arburst[4]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init5 bram5 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[5]),
  .s_axi_awvalid(s_axi_awvalid[5]),
  .s_axi_awaddr (s_axi_awaddr [5]),
  .s_axi_wready (s_axi_wready [5]),
  .s_axi_wvalid (s_axi_wvalid [5]),
  .s_axi_wdata  (s_axi_wdata  [5]),
  .s_axi_wstrb  (s_axi_wstrb  [5]),
  .s_axi_wlast  (s_axi_wlast  [5]),
  .s_axi_bready (s_axi_bready [5]),
  .s_axi_bvalid (s_axi_bvalid [5]),
  .s_axi_bresp  (s_axi_bresp  [5]),
  .s_axi_awlen  (s_axi_awlen  [5]),
  .s_axi_awsize (s_axi_awsize [5]),
  .s_axi_awburst(s_axi_awburst[5]),
  .s_axi_arready(s_axi_arready[5]),
  .s_axi_arvalid(s_axi_arvalid[5]),
  .s_axi_araddr (s_axi_araddr [5]),
  .s_axi_rready (s_axi_rready [5]),
  .s_axi_rvalid (s_axi_rvalid [5]),
  .s_axi_rdata  (s_axi_rdata  [5]),
  .s_axi_rlast  (s_axi_rlast  [5]),
  .s_axi_rresp  (s_axi_rresp  [5]),
  .s_axi_arlen  (s_axi_arlen  [5]),
  .s_axi_arsize (s_axi_arsize [5]),
  .s_axi_arburst(s_axi_arburst[5]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init6 bram6 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[6]),
  .s_axi_awvalid(s_axi_awvalid[6]),
  .s_axi_awaddr (s_axi_awaddr [6]),
  .s_axi_wready (s_axi_wready [6]),
  .s_axi_wvalid (s_axi_wvalid [6]),
  .s_axi_wdata  (s_axi_wdata  [6]),
  .s_axi_wstrb  (s_axi_wstrb  [6]),
  .s_axi_wlast  (s_axi_wlast  [6]),
  .s_axi_bready (s_axi_bready [6]),
  .s_axi_bvalid (s_axi_bvalid [6]),
  .s_axi_bresp  (s_axi_bresp  [6]),
  .s_axi_awlen  (s_axi_awlen  [6]),
  .s_axi_awsize (s_axi_awsize [6]),
  .s_axi_awburst(s_axi_awburst[6]),
  .s_axi_arready(s_axi_arready[6]),
  .s_axi_arvalid(s_axi_arvalid[6]),
  .s_axi_araddr (s_axi_araddr [6]),
  .s_axi_rready (s_axi_rready [6]),
  .s_axi_rvalid (s_axi_rvalid [6]),
  .s_axi_rdata  (s_axi_rdata  [6]),
  .s_axi_rlast  (s_axi_rlast  [6]),
  .s_axi_rresp  (s_axi_rresp  [6]),
  .s_axi_arlen  (s_axi_arlen  [6]),
  .s_axi_arsize (s_axi_arsize [6]),
  .s_axi_arburst(s_axi_arburst[6]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init7 bram7 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[7]),
  .s_axi_awvalid(s_axi_awvalid[7]),
  .s_axi_awaddr (s_axi_awaddr [7]),
  .s_axi_wready (s_axi_wready [7]),
  .s_axi_wvalid (s_axi_wvalid [7]),
  .s_axi_wdata  (s_axi_wdata  [7]),
  .s_axi_wstrb  (s_axi_wstrb  [7]),
  .s_axi_wlast  (s_axi_wlast  [7]),
  .s_axi_bready (s_axi_bready [7]),
  .s_axi_bvalid (s_axi_bvalid [7]),
  .s_axi_bresp  (s_axi_bresp  [7]),
  .s_axi_awlen  (s_axi_awlen  [7]),
  .s_axi_awsize (s_axi_awsize [7]),
  .s_axi_awburst(s_axi_awburst[7]),
  .s_axi_arready(s_axi_arready[7]),
  .s_axi_arvalid(s_axi_arvalid[7]),
  .s_axi_araddr (s_axi_araddr [7]),
  .s_axi_rready (s_axi_rready [7]),
  .s_axi_rvalid (s_axi_rvalid [7]),
  .s_axi_rdata  (s_axi_rdata  [7]),
  .s_axi_rlast  (s_axi_rlast  [7]),
  .s_axi_rresp  (s_axi_rresp  [7]),
  .s_axi_arlen  (s_axi_arlen  [7]),
  .s_axi_arsize (s_axi_arsize [7]),
  .s_axi_arburst(s_axi_arburst[7]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init8 bram8 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[8]),
  .s_axi_awvalid(s_axi_awvalid[8]),
  .s_axi_awaddr (s_axi_awaddr [8]),
  .s_axi_wready (s_axi_wready [8]),
  .s_axi_wvalid (s_axi_wvalid [8]),
  .s_axi_wdata  (s_axi_wdata  [8]),
  .s_axi_wstrb  (s_axi_wstrb  [8]),
  .s_axi_wlast  (s_axi_wlast  [8]),
  .s_axi_bready (s_axi_bready [8]),
  .s_axi_bvalid (s_axi_bvalid [8]),
  .s_axi_bresp  (s_axi_bresp  [8]),
  .s_axi_awlen  (s_axi_awlen  [8]),
  .s_axi_awsize (s_axi_awsize [8]),
  .s_axi_awburst(s_axi_awburst[8]),
  .s_axi_arready(s_axi_arready[8]),
  .s_axi_arvalid(s_axi_arvalid[8]),
  .s_axi_araddr (s_axi_araddr [8]),
  .s_axi_rready (s_axi_rready [8]),
  .s_axi_rvalid (s_axi_rvalid [8]),
  .s_axi_rdata  (s_axi_rdata  [8]),
  .s_axi_rlast  (s_axi_rlast  [8]),
  .s_axi_rresp  (s_axi_rresp  [8]),
  .s_axi_arlen  (s_axi_arlen  [8]),
  .s_axi_arsize (s_axi_arsize [8]),
  .s_axi_arburst(s_axi_arburst[8]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init9 bram9 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[9]),
  .s_axi_awvalid(s_axi_awvalid[9]),
  .s_axi_awaddr (s_axi_awaddr [9]),
  .s_axi_wready (s_axi_wready [9]),
  .s_axi_wvalid (s_axi_wvalid [9]),
  .s_axi_wdata  (s_axi_wdata  [9]),
  .s_axi_wstrb  (s_axi_wstrb  [9]),
  .s_axi_wlast  (s_axi_wlast  [9]),
  .s_axi_bready (s_axi_bready [9]),
  .s_axi_bvalid (s_axi_bvalid [9]),
  .s_axi_bresp  (s_axi_bresp  [9]),
  .s_axi_awlen  (s_axi_awlen  [9]),
  .s_axi_awsize (s_axi_awsize [9]),
  .s_axi_awburst(s_axi_awburst[9]),
  .s_axi_arready(s_axi_arready[9]),
  .s_axi_arvalid(s_axi_arvalid[9]),
  .s_axi_araddr (s_axi_araddr [9]),
  .s_axi_rready (s_axi_rready [9]),
  .s_axi_rvalid (s_axi_rvalid [9]),
  .s_axi_rdata  (s_axi_rdata  [9]),
  .s_axi_rlast  (s_axi_rlast  [9]),
  .s_axi_rresp  (s_axi_rresp  [9]),
  .s_axi_arlen  (s_axi_arlen  [9]),
  .s_axi_arsize (s_axi_arsize [9]),
  .s_axi_arburst(s_axi_arburst[9]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init10 bram10 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[10]),
  .s_axi_awvalid(s_axi_awvalid[10]),
  .s_axi_awaddr (s_axi_awaddr [10]),
  .s_axi_wready (s_axi_wready [10]),
  .s_axi_wvalid (s_axi_wvalid [10]),
  .s_axi_wdata  (s_axi_wdata  [10]),
  .s_axi_wstrb  (s_axi_wstrb  [10]),
  .s_axi_wlast  (s_axi_wlast  [10]),
  .s_axi_bready (s_axi_bready [10]),
  .s_axi_bvalid (s_axi_bvalid [10]),
  .s_axi_bresp  (s_axi_bresp  [10]),
  .s_axi_awlen  (s_axi_awlen  [10]),
  .s_axi_awsize (s_axi_awsize [10]),
  .s_axi_awburst(s_axi_awburst[10]),
  .s_axi_arready(s_axi_arready[10]),
  .s_axi_arvalid(s_axi_arvalid[10]),
  .s_axi_araddr (s_axi_araddr [10]),
  .s_axi_rready (s_axi_rready [10]),
  .s_axi_rvalid (s_axi_rvalid [10]),
  .s_axi_rdata  (s_axi_rdata  [10]),
  .s_axi_rlast  (s_axi_rlast  [10]),
  .s_axi_rresp  (s_axi_rresp  [10]),
  .s_axi_arlen  (s_axi_arlen  [10]),
  .s_axi_arsize (s_axi_arsize [10]),
  .s_axi_arburst(s_axi_arburst[10]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init11 bram11 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[11]),
  .s_axi_awvalid(s_axi_awvalid[11]),
  .s_axi_awaddr (s_axi_awaddr [11]),
  .s_axi_wready (s_axi_wready [11]),
  .s_axi_wvalid (s_axi_wvalid [11]),
  .s_axi_wdata  (s_axi_wdata  [11]),
  .s_axi_wstrb  (s_axi_wstrb  [11]),
  .s_axi_wlast  (s_axi_wlast  [11]),
  .s_axi_bready (s_axi_bready [11]),
  .s_axi_bvalid (s_axi_bvalid [11]),
  .s_axi_bresp  (s_axi_bresp  [11]),
  .s_axi_awlen  (s_axi_awlen  [11]),
  .s_axi_awsize (s_axi_awsize [11]),
  .s_axi_awburst(s_axi_awburst[11]),
  .s_axi_arready(s_axi_arready[11]),
  .s_axi_arvalid(s_axi_arvalid[11]),
  .s_axi_araddr (s_axi_araddr [11]),
  .s_axi_rready (s_axi_rready [11]),
  .s_axi_rvalid (s_axi_rvalid [11]),
  .s_axi_rdata  (s_axi_rdata  [11]),
  .s_axi_rlast  (s_axi_rlast  [11]),
  .s_axi_rresp  (s_axi_rresp  [11]),
  .s_axi_arlen  (s_axi_arlen  [11]),
  .s_axi_arsize (s_axi_arsize [11]),
  .s_axi_arburst(s_axi_arburst[11]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init12 bram12 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[12]),
  .s_axi_awvalid(s_axi_awvalid[12]),
  .s_axi_awaddr (s_axi_awaddr [12]),
  .s_axi_wready (s_axi_wready [12]),
  .s_axi_wvalid (s_axi_wvalid [12]),
  .s_axi_wdata  (s_axi_wdata  [12]),
  .s_axi_wstrb  (s_axi_wstrb  [12]),
  .s_axi_wlast  (s_axi_wlast  [12]),
  .s_axi_bready (s_axi_bready [12]),
  .s_axi_bvalid (s_axi_bvalid [12]),
  .s_axi_bresp  (s_axi_bresp  [12]),
  .s_axi_awlen  (s_axi_awlen  [12]),
  .s_axi_awsize (s_axi_awsize [12]),
  .s_axi_awburst(s_axi_awburst[12]),
  .s_axi_arready(s_axi_arready[12]),
  .s_axi_arvalid(s_axi_arvalid[12]),
  .s_axi_araddr (s_axi_araddr [12]),
  .s_axi_rready (s_axi_rready [12]),
  .s_axi_rvalid (s_axi_rvalid [12]),
  .s_axi_rdata  (s_axi_rdata  [12]),
  .s_axi_rlast  (s_axi_rlast  [12]),
  .s_axi_rresp  (s_axi_rresp  [12]),
  .s_axi_arlen  (s_axi_arlen  [12]),
  .s_axi_arsize (s_axi_arsize [12]),
  .s_axi_arburst(s_axi_arburst[12]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init13 bram13 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[13]),
  .s_axi_awvalid(s_axi_awvalid[13]),
  .s_axi_awaddr (s_axi_awaddr [13]),
  .s_axi_wready (s_axi_wready [13]),
  .s_axi_wvalid (s_axi_wvalid [13]),
  .s_axi_wdata  (s_axi_wdata  [13]),
  .s_axi_wstrb  (s_axi_wstrb  [13]),
  .s_axi_wlast  (s_axi_wlast  [13]),
  .s_axi_bready (s_axi_bready [13]),
  .s_axi_bvalid (s_axi_bvalid [13]),
  .s_axi_bresp  (s_axi_bresp  [13]),
  .s_axi_awlen  (s_axi_awlen  [13]),
  .s_axi_awsize (s_axi_awsize [13]),
  .s_axi_awburst(s_axi_awburst[13]),
  .s_axi_arready(s_axi_arready[13]),
  .s_axi_arvalid(s_axi_arvalid[13]),
  .s_axi_araddr (s_axi_araddr [13]),
  .s_axi_rready (s_axi_rready [13]),
  .s_axi_rvalid (s_axi_rvalid [13]),
  .s_axi_rdata  (s_axi_rdata  [13]),
  .s_axi_rlast  (s_axi_rlast  [13]),
  .s_axi_rresp  (s_axi_rresp  [13]),
  .s_axi_arlen  (s_axi_arlen  [13]),
  .s_axi_arsize (s_axi_arsize [13]),
  .s_axi_arburst(s_axi_arburst[13]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init14 bram14 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[14]),
  .s_axi_awvalid(s_axi_awvalid[14]),
  .s_axi_awaddr (s_axi_awaddr [14]),
  .s_axi_wready (s_axi_wready [14]),
  .s_axi_wvalid (s_axi_wvalid [14]),
  .s_axi_wdata  (s_axi_wdata  [14]),
  .s_axi_wstrb  (s_axi_wstrb  [14]),
  .s_axi_wlast  (s_axi_wlast  [14]),
  .s_axi_bready (s_axi_bready [14]),
  .s_axi_bvalid (s_axi_bvalid [14]),
  .s_axi_bresp  (s_axi_bresp  [14]),
  .s_axi_awlen  (s_axi_awlen  [14]),
  .s_axi_awsize (s_axi_awsize [14]),
  .s_axi_awburst(s_axi_awburst[14]),
  .s_axi_arready(s_axi_arready[14]),
  .s_axi_arvalid(s_axi_arvalid[14]),
  .s_axi_araddr (s_axi_araddr [14]),
  .s_axi_rready (s_axi_rready [14]),
  .s_axi_rvalid (s_axi_rvalid [14]),
  .s_axi_rdata  (s_axi_rdata  [14]),
  .s_axi_rlast  (s_axi_rlast  [14]),
  .s_axi_rresp  (s_axi_rresp  [14]),
  .s_axi_arlen  (s_axi_arlen  [14]),
  .s_axi_arsize (s_axi_arsize [14]),
  .s_axi_arburst(s_axi_arburst[14]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);

bram_init15 bram15 (
  .s_aclk       (hbm_aclk),
  .s_aresetn    (rst_n),
  .s_axi_awready(s_axi_awready[15]),
  .s_axi_awvalid(s_axi_awvalid[15]),
  .s_axi_awaddr (s_axi_awaddr [15]),
  .s_axi_wready (s_axi_wready [15]),
  .s_axi_wvalid (s_axi_wvalid [15]),
  .s_axi_wdata  (s_axi_wdata  [15]),
  .s_axi_wstrb  (s_axi_wstrb  [15]),
  .s_axi_wlast  (s_axi_wlast  [15]),
  .s_axi_bready (s_axi_bready [15]),
  .s_axi_bvalid (s_axi_bvalid [15]),
  .s_axi_bresp  (s_axi_bresp  [15]),
  .s_axi_awlen  (s_axi_awlen  [15]),
  .s_axi_awsize (s_axi_awsize [15]),
  .s_axi_awburst(s_axi_awburst[15]),
  .s_axi_arready(s_axi_arready[15]),
  .s_axi_arvalid(s_axi_arvalid[15]),
  .s_axi_araddr (s_axi_araddr [15]),
  .s_axi_rready (s_axi_rready [15]),
  .s_axi_rvalid (s_axi_rvalid [15]),
  .s_axi_rdata  (s_axi_rdata  [15]),
  .s_axi_rlast  (s_axi_rlast  [15]),
  .s_axi_rresp  (s_axi_rresp  [15]),
  .s_axi_arlen  (s_axi_arlen  [15]),
  .s_axi_arsize (s_axi_arsize [15]),
  .s_axi_arburst(s_axi_arburst[15]),
  .s_axi_awid   (4'd0),
  .s_axi_bid    (),
  .s_axi_arid   (4'd0),
  .s_axi_rid    ()
);
`endif

wire [NUM_GROUP-1:0] launch;
wire [NUM_GROUP-1:0] start_load;
inte #(
  .NUM_GROUP(NUM_GROUP)
) inte_i (
  .sclk          (sclk),
  .xdma_rstn     (xdma_rstn),
  .gpio          (gpio),
  .start_load    (start_load),
  .rst_n         (rst_n),
  .launch        (launch),
  .start_load_all(start_load_all)
);

generate for (genvar m=0; m<NUM_GROUP; m=m+1) begin
  axi_itct axi_itct_i(
    .INTERCONNECT_ACLK   (sclk),
    .INTERCONNECT_ARESETN(rst_n),
    .S00_AXI_ACLK        (sclk),
    .S00_AXI_ARESET_OUT_N(),
    .M00_AXI_ACLK        (hbm_aclk),
    .M00_AXI_ARESET_OUT_N(),
    .S00_AXI_AWREADY     (m_axi_awready[m]),
    .S00_AXI_AWVALID     (m_axi_awvalid[m]),
    .S00_AXI_AWADDR      (m_axi_awaddr [m]),
    .S00_AXI_WREADY      (m_axi_wready [m]),
    .S00_AXI_WVALID      (m_axi_wvalid [m]),
    .S00_AXI_WDATA       (m_axi_wdata  [m]),
    .S00_AXI_WSTRB       (m_axi_wstrb  [m]),
    .S00_AXI_WLAST       (m_axi_wlast  [m]),
    .S00_AXI_BREADY      (m_axi_bready [m]),
    .S00_AXI_BVALID      (m_axi_bvalid [m]),
    .S00_AXI_BRESP       (m_axi_bresp  [m]),
    .S00_AXI_AWLEN       (m_axi_awlen  [m]),
    .S00_AXI_AWSIZE      (m_axi_awsize [m]),
    .S00_AXI_AWBURST     (m_axi_awburst[m]),
    .S00_AXI_AWCACHE     (m_axi_awcache[m]),
    .S00_AXI_ARREADY     (m_axi_arready[m]),
    .S00_AXI_ARVALID     (m_axi_arvalid[m]),
    .S00_AXI_ARADDR      (m_axi_araddr [m]),
    .S00_AXI_RREADY      (m_axi_rready [m]),
    .S00_AXI_RVALID      (m_axi_rvalid [m]),
    .S00_AXI_RDATA       (m_axi_rdata  [m]),
    .S00_AXI_RLAST       (m_axi_rlast  [m]),
    .S00_AXI_RRESP       (m_axi_rresp  [m]),
    .S00_AXI_ARLEN       (m_axi_arlen  [m]),
    .S00_AXI_ARSIZE      (m_axi_arsize [m]),
    .S00_AXI_ARBURST     (m_axi_arburst[m]),
    .S00_AXI_ARCACHE     (m_axi_arcache[m]),
    .S00_AXI_AWID        (1'b0),
    .S00_AXI_BID         (),
    .S00_AXI_AWLOCK      (1'b0),
    .S00_AXI_AWPROT      (3'd0),
    .S00_AXI_AWQOS       (4'd0),
    .S00_AXI_ARID        (1'b0),
    .S00_AXI_RID         (),
    .S00_AXI_ARLOCK      (1'b0),
    .S00_AXI_ARPROT      (3'd0),
    .S00_AXI_ARQOS       (4'd0),
    .M00_AXI_AWREADY     (s_axi_awready[m]),
    .M00_AXI_AWVALID     (s_axi_awvalid[m]),
    .M00_AXI_AWADDR      (s_axi_awaddr [m]),
    .M00_AXI_WREADY      (s_axi_wready [m]),
    .M00_AXI_WVALID      (s_axi_wvalid [m]),
    .M00_AXI_WDATA       (s_axi_wdata  [m]),
    .M00_AXI_WSTRB       (s_axi_wstrb  [m]),
    .M00_AXI_WLAST       (s_axi_wlast  [m]),
    .M00_AXI_BREADY      (s_axi_bready [m]),
    .M00_AXI_BVALID      (s_axi_bvalid [m]),
    .M00_AXI_BRESP       (s_axi_bresp  [m]),
    .M00_AXI_AWLEN       (s_axi_awlen  [m]),
    .M00_AXI_AWSIZE      (s_axi_awsize [m]),
    .M00_AXI_AWBURST     (s_axi_awburst[m]),
    .M00_AXI_AWCACHE     (s_axi_awcache[m]),
    .M00_AXI_ARREADY     (s_axi_arready[m]),
    .M00_AXI_ARVALID     (s_axi_arvalid[m]),
    .M00_AXI_ARADDR      (s_axi_araddr [m]),
    .M00_AXI_RREADY      (s_axi_rready [m]),
    .M00_AXI_RVALID      (s_axi_rvalid [m]),
    .M00_AXI_RDATA       (s_axi_rdata  [m]),
    .M00_AXI_RLAST       (s_axi_rlast  [m]),
    .M00_AXI_RRESP       (s_axi_rresp  [m]),
    .M00_AXI_ARLEN       (s_axi_arlen  [m]),
    .M00_AXI_ARSIZE      (s_axi_arsize [m]),
    .M00_AXI_ARBURST     (s_axi_arburst[m]),
    .M00_AXI_ARCACHE     (s_axi_arcache[m]),
    .M00_AXI_BID         (3'd0),
    .M00_AXI_AWLOCK      (),
    .M00_AXI_AWPROT      (),
    .M00_AXI_AWQOS       (),
    .M00_AXI_AWID        (),
    .M00_AXI_RID         (3'd0),
    .M00_AXI_ARLOCK      (),
    .M00_AXI_ARPROT      (),
    .M00_AXI_ARQOS       (),
    .M00_AXI_ARID        ()
  );
end
endgenerate

/**************************** 数据加载 ****************************/
wire   [NUM_GROUP-1:0] start_turn;
wire   [NUM_GROUP-1:0] done_upload;
wire   [NUM_GROUP-1:0] upload;
wire  [SIZE_GROUP-1:0] wea_load   [NUM_GROUP-1:0];
wire [AWIDTH_BRAM-1:0] addra_load [NUM_GROUP-1:0];
wire [AWIDTH_BRAM-1:0] addrb_load [NUM_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] dout_load  [NUM_GROUP-1:0][SIZE_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] din_load   [NUM_GROUP-1:0][SIZE_GROUP-1:0];
assign upload = start_load; 
generate for (genvar m=0; m<NUM_GROUP; m=m+1) begin
  load #(
    .ID_GROUP   (m),
    .LENGTH     (LENGTH),
    .SIZE_LOOP  (SIZE_LOOP),
    .DWIDTH_FFT (DWIDTH_FFT),
    .SIZE_GROUP (SIZE_GROUP),
    .AWIDTH_HBM (AWIDTH_HBM),
    .DWIDTH_LOAD(DWIDTH_LOAD),
    .DWIDTH_BRAM(DWIDTH_BRAM),
    .AWIDTH_BRAM(AWIDTH_BRAM)
  ) load_i (
    .sclk        (sclk),
    .rst_n       (rst_n),
    .launch      (launch[m]),
    .wea_load    (wea_load[m]),
    .addra_load  (addra_load[m]),
    .addrb_load  (addrb_load[m]),
    .start_load  (start_load[m]),
    .upload      (upload[m]),
    .done_upload (done_upload[m]),

    .dout_load0  (dout_load[m][0]),
    .dout_load1  (dout_load[m][1]),
    .dout_load2  (dout_load[m][2]),
    .dout_load3  (dout_load[m][3]),
    .dout_load4  (dout_load[m][4]),
    .dout_load5  (dout_load[m][5]),
    .dout_load6  (dout_load[m][6]),
    .dout_load7  (dout_load[m][7]),

    .din_load0  (din_load[m][0]),
    .din_load1  (din_load[m][1]),
    .din_load2  (din_load[m][2]),
    .din_load3  (din_load[m][3]),
    .din_load4  (din_load[m][4]),
    .din_load5  (din_load[m][5]),
    .din_load6  (din_load[m][6]),
    .din_load7  (din_load[m][7]),

    .axi_awready(m_axi_awready[m]),
    .axi_awvalid(m_axi_awvalid[m]),
    .axi_awaddr (m_axi_awaddr [m]),
    .axi_awburst(m_axi_awburst[m]),
    .axi_awlen  (m_axi_awlen  [m]),
    .axi_awcache(m_axi_awcache[m]),
    .axi_awsize (m_axi_awsize [m]),
    .axi_wready (m_axi_wready [m]),
    .axi_wvalid (m_axi_wvalid [m]),
    .axi_wdata  (m_axi_wdata  [m]),
    .axi_wstrb  (m_axi_wstrb  [m]),
    .axi_wlast  (m_axi_wlast  [m]),
    .axi_bready (m_axi_bready [m]),
    .axi_bvalid (m_axi_bvalid [m]),
    .axi_bresp  (m_axi_bresp  [m]),
    .axi_arready(m_axi_arready[m]),
    .axi_arvalid(m_axi_arvalid[m]),
    .axi_araddr (m_axi_araddr [m]),
    .axi_arburst(m_axi_arburst[m]),
    .axi_arlen  (m_axi_arlen  [m]),
    .axi_arcache(m_axi_arcache[m]),
    .axi_arsize (m_axi_arsize [m]),
    .axi_rready (m_axi_rready [m]),
    .axi_rvalid (m_axi_rvalid [m]),
    .axi_rdata  (m_axi_rdata  [m]),
    .axi_rlast  (m_axi_rlast  [m]),
    .axi_rresp  (m_axi_rresp  [m])
  );
end
endgenerate

/**************************** 数据缓存 ****************************/
wire   [NUM_GROUP-1:0] web_sw ;
wire [AWIDTH_BRAM-1:0] addrb_sw  [NUM_GROUP-1:0];
wire [AWIDTH_BRAM-1:0] addrb_fft [NUM_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] din_fft   [NUM_GROUP-1:0][SIZE_GROUP-1:0];
wire [DWIDTH_BRAM-1:0] dout_sw   [NUM_GROUP-1:0][SIZE_GROUP-1:0];
generate for (genvar m=0; m<NUM_GROUP; m=m+1) begin
mem #(
  .ID_GROUP   (m),
  .LENGTH     (LENGTH),
  .SIZE_LOOP  (SIZE_LOOP),
  .SIZE_GROUP (SIZE_GROUP),
  .DWIDTH_BRAM(DWIDTH_BRAM),
  .AWIDTH_BRAM(AWIDTH_BRAM)
) mem_i (
  .sclk   (sclk),
  .rst_n  (rst_n),
  .flag0  (1'b0),
  .flag1  (1'b0),

  .wea    (wea_load[m]),
  .addra  (addra_load[m]),
  .dina0  (dout_load[m][0]),
  .dina1  (dout_load[m][1]),
  .dina2  (dout_load[m][2]),
  .dina3  (dout_load[m][3]),
  .dina4  (dout_load[m][4]),
  .dina5  (dout_load[m][5]),
  .dina6  (dout_load[m][6]),
  .dina7  (dout_load[m][7]),

  .web    (web_sw[m]),
  .addrb  (addrb_sw[m]),
  .dinb0  (dout_sw[m][0]),
  .dinb1  (dout_sw[m][1]),
  .dinb2  (dout_sw[m][2]),
  .dinb3  (dout_sw[m][3]),
  .dinb4  (dout_sw[m][4]),
  .dinb5  (dout_sw[m][5]),
  .dinb6  (dout_sw[m][6]),
  .dinb7  (dout_sw[m][7]),

  .addrc  (addrb_load[m]),
  .douta0 (din_load[m][0]),
  .douta1 (din_load[m][1]),
  .douta2 (din_load[m][2]),
  .douta3 (din_load[m][3]),
  .douta4 (din_load[m][4]),
  .douta5 (din_load[m][5]),
  .douta6 (din_load[m][6]),
  .douta7 (din_load[m][7]),

  .addrd  (addrb_fft[m]),
  .doutb0 (din_fft[m][0]),
  .doutb1 (din_fft[m][1]),
  .doutb2 (din_fft[m][2]),
  .doutb3 (din_fft[m][3]),
  .doutb4 (din_fft[m][4]),
  .doutb5 (din_fft[m][5]),
  .doutb6 (din_fft[m][6]),
  .doutb7 (din_fft[m][7])
);
end
endgenerate

/**************************** 数据监控 ****************************/
ila ila_i (
  .clk(sclk),
  .probe0 (m_axi_awready[0]),
  .probe1 (m_axi_awvalid[0]),
  .probe2 (m_axi_awaddr [0]),
  .probe3 (m_axi_wready [0]),
  .probe4 (m_axi_wvalid [0]),
  .probe5 (m_axi_wdata  [0]),
  .probe6 (m_axi_wstrb  [0]),
  .probe7 (m_axi_wlast  [0]),
  .probe8 (m_axi_arready[0]),
  .probe9 (m_axi_arvalid[0]),
  .probe10(m_axi_araddr [0]),
  .probe11(m_axi_rready [0]),
  .probe12(m_axi_rvalid [0]),
  .probe13(m_axi_rdata  [0]),
  .probe14(m_axi_rlast  [0]),
  .probe15(m_axi_awready[15]),
  .probe16(m_axi_awvalid[15]),
  .probe17(m_axi_awaddr [15]),
  .probe18(m_axi_wready [15]),
  .probe19(m_axi_wvalid [15]),
  .probe20(m_axi_wdata  [15]),
  .probe21(m_axi_wstrb  [15]),
  .probe22(m_axi_wlast  [15]),
  .probe23(m_axi_arready[15]),
  .probe24(m_axi_arvalid[15]),
  .probe25(m_axi_araddr [15]),
  .probe26(m_axi_rready [15]),
  .probe27(m_axi_rvalid [15]),
  .probe28(m_axi_rdata  [15]),
  .probe29(m_axi_rlast  [15]),
  .probe30(launch           )
);

endmodule